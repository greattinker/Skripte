// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16;

output N6393,N6402,N6411,N6413,N6322,N6410,N6415,N6407,N6409,N6416;

and AND4 (N17, N15, N3, N6, N5);
nand NAND3 (N18, N17, N1, N10);
nor NOR3 (N19, N15, N9, N16);
nand NAND3 (N20, N1, N8, N6);
and AND2 (N21, N13, N15);
or OR3 (N22, N2, N18, N12);
buf BUF1 (N23, N15);
nand NAND3 (N24, N4, N6, N6);
not NOT1 (N25, N5);
xor XOR2 (N26, N21, N19);
nor NOR2 (N27, N11, N15);
nand NAND2 (N28, N15, N4);
and AND3 (N29, N3, N3, N1);
not NOT1 (N30, N17);
buf BUF1 (N31, N26);
buf BUF1 (N32, N24);
xor XOR2 (N33, N31, N26);
not NOT1 (N34, N27);
nor NOR2 (N35, N22, N15);
or OR3 (N36, N23, N20, N3);
nand NAND2 (N37, N1, N1);
buf BUF1 (N38, N28);
buf BUF1 (N39, N36);
xor XOR2 (N40, N39, N17);
or OR3 (N41, N29, N40, N12);
nand NAND4 (N42, N40, N8, N24, N30);
not NOT1 (N43, N18);
nor NOR3 (N44, N38, N22, N40);
and AND3 (N45, N44, N35, N17);
xor XOR2 (N46, N38, N32);
or OR2 (N47, N29, N45);
xor XOR2 (N48, N43, N5);
not NOT1 (N49, N34);
nor NOR4 (N50, N14, N6, N49, N13);
nor NOR2 (N51, N35, N22);
or OR2 (N52, N50, N28);
not NOT1 (N53, N41);
nor NOR2 (N54, N25, N31);
and AND2 (N55, N47, N42);
xor XOR2 (N56, N5, N27);
not NOT1 (N57, N52);
buf BUF1 (N58, N33);
or OR2 (N59, N56, N8);
or OR4 (N60, N59, N5, N44, N16);
or OR2 (N61, N46, N33);
and AND2 (N62, N48, N17);
nand NAND2 (N63, N57, N55);
nand NAND3 (N64, N6, N23, N55);
buf BUF1 (N65, N51);
buf BUF1 (N66, N62);
buf BUF1 (N67, N54);
not NOT1 (N68, N37);
nor NOR2 (N69, N67, N36);
and AND4 (N70, N64, N26, N34, N58);
not NOT1 (N71, N3);
buf BUF1 (N72, N70);
and AND2 (N73, N65, N13);
not NOT1 (N74, N69);
nand NAND4 (N75, N73, N23, N49, N35);
nand NAND3 (N76, N68, N69, N32);
buf BUF1 (N77, N53);
buf BUF1 (N78, N71);
or OR2 (N79, N66, N14);
nor NOR2 (N80, N79, N16);
buf BUF1 (N81, N61);
not NOT1 (N82, N77);
nand NAND2 (N83, N60, N63);
xor XOR2 (N84, N80, N38);
nor NOR4 (N85, N26, N54, N69, N17);
and AND2 (N86, N81, N13);
xor XOR2 (N87, N78, N53);
or OR4 (N88, N87, N7, N54, N38);
nor NOR2 (N89, N88, N73);
nor NOR4 (N90, N84, N19, N4, N47);
or OR4 (N91, N83, N31, N89, N63);
nand NAND4 (N92, N78, N32, N70, N58);
not NOT1 (N93, N91);
nor NOR4 (N94, N76, N29, N47, N85);
nand NAND4 (N95, N74, N68, N81, N79);
nand NAND3 (N96, N65, N31, N84);
and AND2 (N97, N96, N20);
nor NOR2 (N98, N82, N5);
xor XOR2 (N99, N90, N82);
and AND3 (N100, N97, N6, N40);
nand NAND4 (N101, N92, N22, N54, N55);
xor XOR2 (N102, N94, N47);
nand NAND4 (N103, N86, N101, N86, N86);
not NOT1 (N104, N51);
and AND4 (N105, N102, N73, N103, N27);
nor NOR3 (N106, N1, N58, N35);
nand NAND4 (N107, N93, N70, N32, N43);
buf BUF1 (N108, N98);
xor XOR2 (N109, N95, N81);
xor XOR2 (N110, N100, N26);
nor NOR3 (N111, N106, N26, N9);
nor NOR3 (N112, N110, N105, N80);
and AND4 (N113, N54, N50, N47, N39);
or OR4 (N114, N108, N17, N63, N32);
or OR2 (N115, N99, N14);
xor XOR2 (N116, N75, N11);
not NOT1 (N117, N104);
and AND2 (N118, N109, N49);
xor XOR2 (N119, N114, N96);
or OR2 (N120, N115, N118);
and AND3 (N121, N115, N61, N98);
nand NAND3 (N122, N117, N12, N43);
or OR3 (N123, N107, N52, N62);
nor NOR3 (N124, N122, N2, N7);
buf BUF1 (N125, N123);
nor NOR2 (N126, N119, N101);
not NOT1 (N127, N112);
buf BUF1 (N128, N111);
or OR2 (N129, N124, N33);
and AND4 (N130, N126, N78, N95, N3);
nor NOR3 (N131, N127, N123, N79);
or OR3 (N132, N121, N87, N81);
and AND4 (N133, N72, N26, N57, N78);
buf BUF1 (N134, N131);
nand NAND3 (N135, N128, N125, N102);
not NOT1 (N136, N102);
nand NAND3 (N137, N136, N133, N52);
nand NAND4 (N138, N28, N63, N85, N96);
buf BUF1 (N139, N137);
or OR4 (N140, N129, N70, N94, N43);
nor NOR2 (N141, N134, N107);
nand NAND4 (N142, N135, N129, N77, N118);
buf BUF1 (N143, N140);
nor NOR3 (N144, N142, N140, N62);
xor XOR2 (N145, N120, N107);
or OR3 (N146, N116, N50, N96);
xor XOR2 (N147, N143, N50);
not NOT1 (N148, N141);
nor NOR4 (N149, N138, N114, N2, N91);
xor XOR2 (N150, N147, N102);
buf BUF1 (N151, N113);
and AND4 (N152, N130, N142, N50, N46);
not NOT1 (N153, N144);
or OR2 (N154, N151, N1);
buf BUF1 (N155, N149);
nand NAND4 (N156, N150, N3, N35, N94);
and AND2 (N157, N156, N41);
not NOT1 (N158, N132);
and AND4 (N159, N145, N7, N114, N147);
or OR4 (N160, N158, N79, N135, N142);
or OR3 (N161, N155, N151, N82);
nand NAND2 (N162, N146, N22);
xor XOR2 (N163, N154, N33);
buf BUF1 (N164, N162);
nand NAND3 (N165, N152, N95, N32);
nor NOR3 (N166, N153, N111, N152);
nand NAND3 (N167, N148, N90, N55);
not NOT1 (N168, N139);
nand NAND2 (N169, N160, N115);
nand NAND4 (N170, N161, N141, N107, N12);
buf BUF1 (N171, N168);
and AND3 (N172, N167, N150, N77);
or OR3 (N173, N165, N167, N19);
xor XOR2 (N174, N171, N16);
and AND4 (N175, N164, N32, N158, N59);
buf BUF1 (N176, N163);
not NOT1 (N177, N166);
buf BUF1 (N178, N172);
nor NOR2 (N179, N157, N18);
xor XOR2 (N180, N175, N25);
or OR2 (N181, N159, N94);
nand NAND2 (N182, N173, N94);
buf BUF1 (N183, N177);
and AND3 (N184, N178, N88, N75);
xor XOR2 (N185, N174, N40);
buf BUF1 (N186, N169);
nor NOR2 (N187, N184, N49);
not NOT1 (N188, N176);
or OR4 (N189, N170, N184, N110, N91);
and AND3 (N190, N183, N182, N43);
nand NAND4 (N191, N136, N131, N121, N51);
buf BUF1 (N192, N190);
or OR2 (N193, N188, N159);
nor NOR2 (N194, N179, N148);
nor NOR2 (N195, N185, N53);
buf BUF1 (N196, N181);
buf BUF1 (N197, N195);
or OR4 (N198, N191, N88, N154, N72);
nor NOR2 (N199, N197, N67);
buf BUF1 (N200, N187);
xor XOR2 (N201, N199, N61);
buf BUF1 (N202, N194);
nor NOR2 (N203, N189, N133);
buf BUF1 (N204, N202);
and AND2 (N205, N200, N119);
nand NAND4 (N206, N193, N101, N156, N44);
buf BUF1 (N207, N203);
not NOT1 (N208, N196);
or OR3 (N209, N207, N117, N43);
buf BUF1 (N210, N201);
and AND3 (N211, N205, N133, N18);
or OR3 (N212, N206, N60, N21);
buf BUF1 (N213, N186);
nor NOR2 (N214, N198, N126);
nand NAND2 (N215, N208, N118);
and AND3 (N216, N215, N213, N179);
or OR2 (N217, N145, N50);
nor NOR3 (N218, N209, N198, N177);
xor XOR2 (N219, N212, N86);
nand NAND2 (N220, N180, N65);
and AND4 (N221, N217, N110, N16, N17);
nor NOR4 (N222, N219, N15, N32, N23);
buf BUF1 (N223, N192);
nand NAND3 (N224, N220, N201, N84);
and AND4 (N225, N224, N57, N194, N5);
buf BUF1 (N226, N210);
and AND4 (N227, N221, N197, N4, N13);
not NOT1 (N228, N223);
xor XOR2 (N229, N214, N137);
buf BUF1 (N230, N226);
or OR4 (N231, N230, N65, N78, N119);
not NOT1 (N232, N218);
not NOT1 (N233, N231);
not NOT1 (N234, N228);
xor XOR2 (N235, N211, N123);
not NOT1 (N236, N233);
buf BUF1 (N237, N225);
not NOT1 (N238, N222);
buf BUF1 (N239, N234);
buf BUF1 (N240, N227);
nand NAND2 (N241, N229, N114);
nand NAND4 (N242, N236, N108, N188, N8);
nand NAND4 (N243, N240, N37, N108, N105);
or OR2 (N244, N238, N45);
buf BUF1 (N245, N239);
nand NAND3 (N246, N241, N175, N208);
nor NOR4 (N247, N245, N182, N33, N213);
nand NAND3 (N248, N232, N2, N22);
buf BUF1 (N249, N243);
nor NOR2 (N250, N248, N174);
xor XOR2 (N251, N249, N204);
or OR3 (N252, N20, N2, N95);
xor XOR2 (N253, N246, N8);
and AND4 (N254, N216, N80, N14, N161);
nor NOR4 (N255, N247, N193, N148, N196);
or OR2 (N256, N250, N72);
nor NOR3 (N257, N235, N86, N20);
nand NAND2 (N258, N237, N43);
nor NOR4 (N259, N257, N12, N126, N77);
or OR4 (N260, N256, N212, N1, N202);
nor NOR3 (N261, N253, N163, N119);
not NOT1 (N262, N254);
not NOT1 (N263, N252);
nand NAND3 (N264, N258, N186, N27);
buf BUF1 (N265, N260);
or OR2 (N266, N264, N191);
and AND4 (N267, N261, N239, N194, N159);
xor XOR2 (N268, N251, N148);
or OR3 (N269, N263, N50, N167);
not NOT1 (N270, N244);
or OR4 (N271, N266, N73, N202, N37);
xor XOR2 (N272, N269, N77);
and AND4 (N273, N272, N159, N139, N112);
and AND3 (N274, N255, N115, N180);
not NOT1 (N275, N273);
not NOT1 (N276, N270);
and AND2 (N277, N242, N146);
buf BUF1 (N278, N268);
buf BUF1 (N279, N271);
and AND4 (N280, N277, N81, N119, N58);
nor NOR4 (N281, N259, N119, N278, N99);
not NOT1 (N282, N44);
or OR3 (N283, N281, N3, N172);
nand NAND3 (N284, N275, N254, N155);
buf BUF1 (N285, N284);
and AND4 (N286, N279, N203, N201, N83);
xor XOR2 (N287, N286, N172);
and AND2 (N288, N265, N84);
xor XOR2 (N289, N285, N169);
not NOT1 (N290, N276);
or OR3 (N291, N280, N34, N253);
buf BUF1 (N292, N274);
and AND2 (N293, N267, N187);
buf BUF1 (N294, N290);
not NOT1 (N295, N287);
and AND4 (N296, N291, N189, N240, N131);
xor XOR2 (N297, N289, N175);
and AND3 (N298, N296, N77, N222);
and AND3 (N299, N297, N268, N51);
xor XOR2 (N300, N294, N264);
or OR2 (N301, N299, N208);
buf BUF1 (N302, N298);
xor XOR2 (N303, N300, N192);
nor NOR2 (N304, N288, N192);
not NOT1 (N305, N292);
not NOT1 (N306, N283);
or OR2 (N307, N262, N127);
xor XOR2 (N308, N305, N39);
or OR3 (N309, N303, N113, N213);
xor XOR2 (N310, N306, N253);
xor XOR2 (N311, N310, N93);
or OR3 (N312, N308, N134, N227);
xor XOR2 (N313, N301, N124);
or OR3 (N314, N293, N35, N245);
xor XOR2 (N315, N313, N105);
not NOT1 (N316, N302);
not NOT1 (N317, N311);
or OR4 (N318, N309, N253, N161, N217);
nor NOR2 (N319, N295, N102);
buf BUF1 (N320, N282);
or OR2 (N321, N317, N66);
nor NOR3 (N322, N315, N105, N247);
and AND4 (N323, N314, N291, N2, N65);
nor NOR2 (N324, N320, N203);
buf BUF1 (N325, N316);
buf BUF1 (N326, N318);
nand NAND2 (N327, N319, N227);
not NOT1 (N328, N324);
xor XOR2 (N329, N323, N280);
not NOT1 (N330, N325);
nand NAND2 (N331, N304, N222);
xor XOR2 (N332, N312, N309);
nand NAND2 (N333, N329, N154);
not NOT1 (N334, N307);
nand NAND3 (N335, N322, N297, N176);
xor XOR2 (N336, N321, N201);
or OR2 (N337, N336, N118);
not NOT1 (N338, N330);
nand NAND4 (N339, N327, N269, N102, N82);
nor NOR4 (N340, N338, N208, N56, N54);
not NOT1 (N341, N326);
or OR2 (N342, N335, N293);
not NOT1 (N343, N328);
buf BUF1 (N344, N337);
nand NAND2 (N345, N341, N339);
xor XOR2 (N346, N102, N204);
xor XOR2 (N347, N346, N144);
nand NAND3 (N348, N333, N266, N79);
buf BUF1 (N349, N334);
and AND3 (N350, N349, N323, N113);
buf BUF1 (N351, N347);
or OR3 (N352, N340, N2, N206);
not NOT1 (N353, N351);
nor NOR4 (N354, N345, N122, N230, N14);
xor XOR2 (N355, N343, N12);
buf BUF1 (N356, N355);
nor NOR4 (N357, N344, N32, N92, N35);
and AND3 (N358, N348, N305, N270);
and AND4 (N359, N342, N294, N203, N317);
nand NAND3 (N360, N352, N49, N178);
or OR3 (N361, N357, N114, N85);
nor NOR3 (N362, N331, N85, N23);
or OR4 (N363, N353, N303, N218, N219);
and AND4 (N364, N356, N251, N176, N308);
not NOT1 (N365, N358);
and AND4 (N366, N363, N256, N101, N76);
xor XOR2 (N367, N366, N225);
or OR2 (N368, N359, N334);
xor XOR2 (N369, N332, N122);
nor NOR4 (N370, N361, N73, N50, N210);
xor XOR2 (N371, N365, N25);
and AND4 (N372, N371, N131, N294, N257);
nand NAND3 (N373, N360, N366, N97);
nor NOR3 (N374, N370, N250, N342);
buf BUF1 (N375, N373);
xor XOR2 (N376, N375, N298);
and AND2 (N377, N362, N67);
not NOT1 (N378, N367);
buf BUF1 (N379, N368);
not NOT1 (N380, N379);
nor NOR2 (N381, N376, N30);
xor XOR2 (N382, N369, N280);
xor XOR2 (N383, N372, N267);
nand NAND2 (N384, N364, N265);
xor XOR2 (N385, N382, N368);
or OR3 (N386, N378, N108, N117);
xor XOR2 (N387, N386, N61);
nor NOR2 (N388, N354, N249);
not NOT1 (N389, N381);
nand NAND4 (N390, N385, N363, N369, N179);
nor NOR4 (N391, N374, N4, N202, N195);
and AND4 (N392, N387, N85, N25, N328);
xor XOR2 (N393, N384, N382);
or OR4 (N394, N390, N320, N46, N33);
buf BUF1 (N395, N391);
and AND2 (N396, N393, N66);
not NOT1 (N397, N380);
xor XOR2 (N398, N394, N73);
not NOT1 (N399, N383);
not NOT1 (N400, N399);
and AND4 (N401, N350, N312, N209, N69);
and AND2 (N402, N396, N320);
nand NAND2 (N403, N395, N227);
and AND3 (N404, N400, N336, N8);
and AND2 (N405, N388, N398);
or OR4 (N406, N167, N1, N293, N22);
not NOT1 (N407, N405);
nor NOR4 (N408, N389, N295, N90, N248);
and AND2 (N409, N402, N327);
nand NAND4 (N410, N377, N357, N159, N292);
xor XOR2 (N411, N392, N384);
nor NOR2 (N412, N404, N198);
or OR3 (N413, N406, N21, N281);
not NOT1 (N414, N401);
not NOT1 (N415, N408);
nor NOR3 (N416, N407, N152, N374);
or OR3 (N417, N410, N372, N27);
and AND2 (N418, N403, N220);
xor XOR2 (N419, N411, N142);
and AND4 (N420, N418, N88, N413, N57);
nand NAND3 (N421, N325, N36, N400);
not NOT1 (N422, N420);
nor NOR3 (N423, N416, N361, N406);
or OR2 (N424, N415, N327);
xor XOR2 (N425, N419, N248);
xor XOR2 (N426, N417, N87);
or OR4 (N427, N409, N298, N393, N258);
nand NAND2 (N428, N414, N348);
nand NAND4 (N429, N426, N94, N382, N15);
not NOT1 (N430, N421);
nor NOR2 (N431, N424, N120);
buf BUF1 (N432, N423);
xor XOR2 (N433, N425, N354);
buf BUF1 (N434, N422);
nor NOR3 (N435, N427, N189, N1);
xor XOR2 (N436, N412, N301);
and AND2 (N437, N434, N356);
and AND3 (N438, N430, N64, N91);
nand NAND4 (N439, N431, N308, N379, N101);
nor NOR4 (N440, N438, N86, N99, N395);
buf BUF1 (N441, N433);
or OR3 (N442, N439, N380, N3);
nor NOR3 (N443, N397, N326, N245);
nand NAND3 (N444, N435, N194, N371);
or OR4 (N445, N432, N334, N240, N387);
xor XOR2 (N446, N428, N88);
xor XOR2 (N447, N445, N217);
and AND3 (N448, N447, N130, N4);
and AND3 (N449, N443, N178, N399);
buf BUF1 (N450, N436);
nand NAND4 (N451, N441, N221, N33, N214);
and AND4 (N452, N448, N404, N438, N165);
buf BUF1 (N453, N449);
and AND2 (N454, N450, N275);
xor XOR2 (N455, N444, N81);
and AND4 (N456, N454, N125, N211, N89);
or OR4 (N457, N446, N418, N392, N389);
xor XOR2 (N458, N429, N388);
or OR4 (N459, N456, N321, N345, N218);
xor XOR2 (N460, N452, N239);
xor XOR2 (N461, N451, N367);
buf BUF1 (N462, N461);
xor XOR2 (N463, N458, N290);
nor NOR3 (N464, N457, N179, N400);
not NOT1 (N465, N440);
buf BUF1 (N466, N442);
and AND4 (N467, N464, N200, N47, N221);
xor XOR2 (N468, N466, N393);
and AND3 (N469, N463, N61, N87);
nand NAND2 (N470, N468, N414);
nor NOR4 (N471, N462, N238, N109, N370);
buf BUF1 (N472, N471);
nand NAND2 (N473, N437, N254);
not NOT1 (N474, N470);
xor XOR2 (N475, N455, N225);
buf BUF1 (N476, N472);
nand NAND2 (N477, N473, N102);
and AND2 (N478, N475, N141);
buf BUF1 (N479, N474);
nand NAND3 (N480, N479, N3, N184);
buf BUF1 (N481, N453);
nand NAND4 (N482, N467, N335, N87, N319);
nor NOR3 (N483, N476, N269, N7);
not NOT1 (N484, N477);
and AND4 (N485, N459, N131, N144, N136);
or OR2 (N486, N480, N434);
or OR3 (N487, N485, N431, N234);
or OR3 (N488, N465, N455, N374);
not NOT1 (N489, N482);
or OR2 (N490, N486, N98);
nand NAND2 (N491, N484, N462);
nand NAND2 (N492, N487, N65);
and AND4 (N493, N460, N245, N49, N245);
or OR2 (N494, N488, N14);
and AND4 (N495, N491, N228, N340, N38);
nor NOR4 (N496, N481, N295, N144, N378);
xor XOR2 (N497, N489, N104);
and AND3 (N498, N495, N493, N295);
nand NAND4 (N499, N379, N259, N281, N485);
xor XOR2 (N500, N483, N412);
or OR3 (N501, N469, N207, N136);
buf BUF1 (N502, N501);
xor XOR2 (N503, N497, N258);
and AND4 (N504, N478, N96, N497, N159);
xor XOR2 (N505, N496, N472);
or OR4 (N506, N503, N284, N318, N240);
xor XOR2 (N507, N490, N474);
nor NOR3 (N508, N492, N161, N456);
or OR3 (N509, N508, N314, N69);
and AND2 (N510, N494, N144);
or OR3 (N511, N509, N485, N289);
nand NAND4 (N512, N504, N115, N227, N166);
xor XOR2 (N513, N502, N256);
buf BUF1 (N514, N498);
buf BUF1 (N515, N512);
buf BUF1 (N516, N515);
xor XOR2 (N517, N511, N341);
buf BUF1 (N518, N505);
and AND2 (N519, N499, N516);
nor NOR2 (N520, N301, N8);
not NOT1 (N521, N507);
or OR2 (N522, N519, N262);
xor XOR2 (N523, N510, N363);
xor XOR2 (N524, N500, N482);
buf BUF1 (N525, N523);
xor XOR2 (N526, N518, N111);
nor NOR2 (N527, N524, N69);
and AND2 (N528, N517, N87);
xor XOR2 (N529, N506, N518);
and AND4 (N530, N526, N249, N401, N206);
and AND3 (N531, N520, N83, N196);
not NOT1 (N532, N527);
nand NAND2 (N533, N531, N332);
and AND3 (N534, N525, N171, N230);
and AND2 (N535, N529, N126);
or OR4 (N536, N532, N135, N148, N355);
not NOT1 (N537, N535);
not NOT1 (N538, N522);
nor NOR4 (N539, N534, N17, N433, N241);
and AND4 (N540, N528, N316, N495, N193);
not NOT1 (N541, N540);
not NOT1 (N542, N533);
and AND4 (N543, N541, N102, N257, N435);
nor NOR2 (N544, N514, N23);
or OR3 (N545, N543, N194, N402);
xor XOR2 (N546, N521, N539);
nor NOR4 (N547, N458, N330, N339, N356);
not NOT1 (N548, N542);
buf BUF1 (N549, N547);
nor NOR3 (N550, N549, N490, N414);
and AND2 (N551, N550, N198);
nor NOR2 (N552, N537, N52);
or OR2 (N553, N545, N144);
not NOT1 (N554, N551);
not NOT1 (N555, N538);
buf BUF1 (N556, N536);
nor NOR3 (N557, N530, N195, N491);
not NOT1 (N558, N553);
and AND3 (N559, N513, N10, N195);
or OR2 (N560, N554, N367);
and AND4 (N561, N544, N545, N408, N514);
not NOT1 (N562, N546);
buf BUF1 (N563, N555);
xor XOR2 (N564, N556, N247);
nor NOR2 (N565, N557, N350);
and AND3 (N566, N562, N177, N260);
xor XOR2 (N567, N561, N118);
not NOT1 (N568, N567);
not NOT1 (N569, N565);
xor XOR2 (N570, N559, N428);
not NOT1 (N571, N548);
xor XOR2 (N572, N568, N302);
not NOT1 (N573, N569);
nor NOR4 (N574, N570, N518, N194, N76);
not NOT1 (N575, N571);
nor NOR2 (N576, N575, N399);
xor XOR2 (N577, N560, N255);
nor NOR4 (N578, N576, N276, N345, N547);
nand NAND4 (N579, N564, N201, N383, N63);
xor XOR2 (N580, N573, N278);
and AND2 (N581, N558, N531);
xor XOR2 (N582, N577, N24);
not NOT1 (N583, N574);
or OR2 (N584, N566, N368);
and AND3 (N585, N572, N550, N150);
not NOT1 (N586, N579);
buf BUF1 (N587, N563);
or OR2 (N588, N587, N509);
nand NAND3 (N589, N586, N80, N327);
or OR2 (N590, N588, N498);
buf BUF1 (N591, N589);
nor NOR3 (N592, N582, N577, N591);
xor XOR2 (N593, N399, N359);
nor NOR4 (N594, N584, N395, N317, N536);
nand NAND2 (N595, N592, N367);
not NOT1 (N596, N583);
buf BUF1 (N597, N580);
or OR3 (N598, N581, N211, N458);
xor XOR2 (N599, N578, N191);
nor NOR2 (N600, N599, N517);
and AND3 (N601, N597, N122, N2);
or OR3 (N602, N552, N180, N246);
and AND3 (N603, N600, N94, N95);
not NOT1 (N604, N590);
nor NOR3 (N605, N602, N216, N82);
not NOT1 (N606, N596);
not NOT1 (N607, N598);
nand NAND3 (N608, N603, N585, N43);
not NOT1 (N609, N527);
xor XOR2 (N610, N607, N555);
or OR2 (N611, N610, N204);
nand NAND2 (N612, N609, N522);
not NOT1 (N613, N604);
xor XOR2 (N614, N606, N479);
nor NOR4 (N615, N613, N598, N378, N79);
xor XOR2 (N616, N594, N520);
nor NOR2 (N617, N612, N355);
and AND3 (N618, N595, N75, N77);
xor XOR2 (N619, N617, N407);
nor NOR2 (N620, N593, N418);
not NOT1 (N621, N616);
not NOT1 (N622, N621);
nor NOR3 (N623, N611, N350, N415);
buf BUF1 (N624, N620);
xor XOR2 (N625, N619, N418);
nor NOR4 (N626, N625, N599, N10, N330);
buf BUF1 (N627, N601);
not NOT1 (N628, N624);
nor NOR3 (N629, N626, N220, N331);
not NOT1 (N630, N608);
or OR4 (N631, N622, N312, N199, N603);
nand NAND3 (N632, N614, N170, N440);
or OR2 (N633, N615, N408);
nand NAND3 (N634, N618, N30, N282);
buf BUF1 (N635, N623);
and AND3 (N636, N605, N118, N539);
nand NAND4 (N637, N636, N607, N531, N139);
and AND2 (N638, N630, N284);
and AND3 (N639, N632, N164, N521);
nor NOR2 (N640, N638, N398);
nand NAND3 (N641, N637, N5, N462);
and AND3 (N642, N628, N109, N484);
buf BUF1 (N643, N639);
and AND2 (N644, N640, N347);
or OR3 (N645, N633, N369, N5);
and AND4 (N646, N631, N555, N117, N428);
or OR3 (N647, N629, N239, N626);
buf BUF1 (N648, N641);
nor NOR4 (N649, N635, N18, N366, N205);
nor NOR2 (N650, N643, N571);
or OR4 (N651, N649, N252, N76, N203);
and AND2 (N652, N650, N171);
or OR3 (N653, N644, N17, N320);
nand NAND4 (N654, N647, N369, N334, N400);
nand NAND4 (N655, N651, N160, N321, N639);
and AND4 (N656, N653, N135, N195, N28);
nand NAND3 (N657, N654, N191, N499);
buf BUF1 (N658, N634);
nor NOR3 (N659, N657, N230, N306);
not NOT1 (N660, N642);
buf BUF1 (N661, N659);
xor XOR2 (N662, N627, N609);
xor XOR2 (N663, N646, N617);
buf BUF1 (N664, N656);
nand NAND2 (N665, N663, N649);
nand NAND2 (N666, N661, N372);
nor NOR3 (N667, N664, N89, N318);
xor XOR2 (N668, N660, N587);
buf BUF1 (N669, N658);
nand NAND4 (N670, N669, N359, N152, N97);
xor XOR2 (N671, N662, N534);
nor NOR3 (N672, N671, N467, N270);
xor XOR2 (N673, N665, N208);
and AND4 (N674, N670, N31, N645, N598);
nand NAND2 (N675, N2, N12);
or OR3 (N676, N675, N505, N151);
or OR2 (N677, N652, N246);
or OR4 (N678, N655, N178, N658, N228);
not NOT1 (N679, N677);
nor NOR3 (N680, N674, N377, N3);
and AND3 (N681, N676, N425, N368);
buf BUF1 (N682, N666);
and AND2 (N683, N682, N295);
and AND3 (N684, N648, N200, N487);
or OR3 (N685, N679, N199, N555);
buf BUF1 (N686, N672);
and AND2 (N687, N686, N151);
xor XOR2 (N688, N678, N602);
and AND2 (N689, N687, N166);
nand NAND3 (N690, N684, N289, N132);
nor NOR3 (N691, N667, N329, N263);
buf BUF1 (N692, N681);
not NOT1 (N693, N690);
and AND4 (N694, N688, N504, N294, N657);
nand NAND2 (N695, N673, N645);
not NOT1 (N696, N694);
buf BUF1 (N697, N695);
nor NOR3 (N698, N683, N278, N33);
not NOT1 (N699, N698);
xor XOR2 (N700, N689, N158);
nor NOR4 (N701, N691, N609, N411, N290);
or OR3 (N702, N692, N564, N32);
or OR4 (N703, N685, N654, N213, N547);
buf BUF1 (N704, N699);
or OR2 (N705, N696, N502);
and AND3 (N706, N703, N238, N67);
and AND4 (N707, N706, N189, N421, N302);
xor XOR2 (N708, N668, N306);
nor NOR4 (N709, N702, N75, N252, N426);
or OR3 (N710, N707, N158, N544);
xor XOR2 (N711, N704, N597);
xor XOR2 (N712, N710, N167);
and AND4 (N713, N711, N39, N672, N76);
and AND4 (N714, N713, N1, N9, N625);
nand NAND3 (N715, N714, N579, N11);
nand NAND3 (N716, N701, N323, N78);
and AND4 (N717, N705, N360, N641, N327);
xor XOR2 (N718, N712, N76);
not NOT1 (N719, N700);
not NOT1 (N720, N693);
not NOT1 (N721, N716);
nand NAND4 (N722, N721, N591, N437, N510);
or OR2 (N723, N717, N331);
and AND3 (N724, N723, N500, N346);
buf BUF1 (N725, N719);
nor NOR2 (N726, N725, N384);
xor XOR2 (N727, N709, N363);
buf BUF1 (N728, N724);
xor XOR2 (N729, N718, N118);
not NOT1 (N730, N728);
nor NOR3 (N731, N730, N118, N709);
nand NAND3 (N732, N731, N68, N128);
xor XOR2 (N733, N697, N332);
and AND3 (N734, N729, N722, N269);
not NOT1 (N735, N139);
buf BUF1 (N736, N735);
or OR4 (N737, N715, N402, N456, N285);
or OR4 (N738, N733, N607, N696, N675);
buf BUF1 (N739, N732);
buf BUF1 (N740, N736);
buf BUF1 (N741, N680);
nand NAND2 (N742, N737, N408);
or OR2 (N743, N727, N401);
and AND2 (N744, N708, N453);
nor NOR3 (N745, N744, N420, N60);
nor NOR2 (N746, N741, N387);
nor NOR4 (N747, N726, N374, N47, N11);
nor NOR4 (N748, N747, N743, N518, N171);
and AND3 (N749, N34, N108, N70);
not NOT1 (N750, N738);
or OR4 (N751, N720, N433, N157, N271);
buf BUF1 (N752, N742);
and AND2 (N753, N749, N565);
buf BUF1 (N754, N750);
nor NOR4 (N755, N745, N133, N98, N685);
and AND4 (N756, N746, N628, N45, N197);
nor NOR4 (N757, N753, N75, N247, N369);
nor NOR2 (N758, N740, N169);
xor XOR2 (N759, N757, N232);
xor XOR2 (N760, N751, N749);
not NOT1 (N761, N734);
buf BUF1 (N762, N758);
or OR2 (N763, N755, N629);
and AND4 (N764, N739, N590, N375, N763);
nor NOR2 (N765, N763, N592);
xor XOR2 (N766, N756, N410);
and AND3 (N767, N754, N43, N647);
xor XOR2 (N768, N752, N606);
buf BUF1 (N769, N761);
or OR2 (N770, N760, N500);
xor XOR2 (N771, N770, N701);
xor XOR2 (N772, N765, N549);
not NOT1 (N773, N772);
or OR2 (N774, N771, N430);
xor XOR2 (N775, N768, N444);
and AND2 (N776, N748, N221);
xor XOR2 (N777, N762, N530);
nor NOR4 (N778, N775, N675, N219, N67);
or OR2 (N779, N773, N74);
or OR3 (N780, N778, N673, N505);
nor NOR2 (N781, N777, N569);
nand NAND3 (N782, N769, N14, N21);
and AND2 (N783, N776, N485);
buf BUF1 (N784, N782);
or OR2 (N785, N781, N706);
nand NAND3 (N786, N783, N16, N742);
buf BUF1 (N787, N774);
nor NOR2 (N788, N759, N628);
nor NOR2 (N789, N764, N181);
and AND3 (N790, N785, N589, N740);
or OR3 (N791, N790, N248, N17);
or OR3 (N792, N788, N711, N470);
nor NOR3 (N793, N792, N625, N116);
xor XOR2 (N794, N779, N191);
nand NAND2 (N795, N784, N324);
nor NOR4 (N796, N794, N665, N408, N611);
xor XOR2 (N797, N766, N675);
xor XOR2 (N798, N793, N13);
nand NAND4 (N799, N795, N17, N449, N87);
or OR4 (N800, N796, N669, N154, N98);
or OR4 (N801, N799, N197, N231, N134);
and AND4 (N802, N767, N579, N228, N392);
not NOT1 (N803, N802);
xor XOR2 (N804, N798, N770);
buf BUF1 (N805, N803);
and AND4 (N806, N801, N561, N93, N597);
and AND4 (N807, N780, N195, N417, N636);
nand NAND3 (N808, N786, N490, N330);
and AND3 (N809, N789, N218, N415);
and AND3 (N810, N800, N166, N586);
or OR2 (N811, N808, N376);
buf BUF1 (N812, N807);
xor XOR2 (N813, N797, N71);
nand NAND2 (N814, N813, N327);
nor NOR3 (N815, N811, N247, N49);
nor NOR3 (N816, N787, N531, N25);
and AND4 (N817, N805, N71, N37, N699);
nand NAND2 (N818, N804, N509);
xor XOR2 (N819, N817, N451);
and AND2 (N820, N814, N317);
nand NAND3 (N821, N812, N101, N526);
buf BUF1 (N822, N816);
nand NAND3 (N823, N820, N135, N144);
nand NAND2 (N824, N810, N609);
nor NOR4 (N825, N822, N110, N570, N782);
and AND4 (N826, N791, N130, N261, N442);
nand NAND4 (N827, N824, N783, N176, N806);
buf BUF1 (N828, N61);
buf BUF1 (N829, N823);
xor XOR2 (N830, N826, N360);
not NOT1 (N831, N830);
xor XOR2 (N832, N829, N661);
xor XOR2 (N833, N827, N145);
and AND2 (N834, N821, N478);
not NOT1 (N835, N819);
nor NOR2 (N836, N832, N685);
xor XOR2 (N837, N833, N495);
nand NAND3 (N838, N834, N433, N81);
nor NOR3 (N839, N815, N694, N157);
and AND2 (N840, N818, N803);
nor NOR3 (N841, N825, N508, N633);
or OR4 (N842, N839, N527, N417, N217);
buf BUF1 (N843, N836);
buf BUF1 (N844, N838);
buf BUF1 (N845, N844);
or OR2 (N846, N837, N153);
xor XOR2 (N847, N831, N532);
nor NOR4 (N848, N828, N579, N273, N733);
and AND2 (N849, N846, N801);
nand NAND4 (N850, N840, N566, N60, N606);
and AND4 (N851, N843, N675, N633, N37);
buf BUF1 (N852, N848);
not NOT1 (N853, N842);
or OR3 (N854, N809, N775, N541);
nand NAND4 (N855, N841, N311, N610, N119);
not NOT1 (N856, N847);
not NOT1 (N857, N854);
xor XOR2 (N858, N855, N841);
or OR4 (N859, N852, N256, N537, N176);
and AND4 (N860, N850, N782, N817, N558);
buf BUF1 (N861, N856);
or OR4 (N862, N861, N564, N634, N194);
buf BUF1 (N863, N859);
and AND4 (N864, N853, N37, N457, N384);
and AND4 (N865, N857, N63, N403, N779);
xor XOR2 (N866, N860, N328);
buf BUF1 (N867, N864);
not NOT1 (N868, N863);
not NOT1 (N869, N858);
not NOT1 (N870, N866);
nand NAND3 (N871, N867, N224, N696);
and AND3 (N872, N851, N737, N262);
nor NOR4 (N873, N862, N212, N444, N117);
buf BUF1 (N874, N873);
and AND3 (N875, N865, N775, N803);
and AND4 (N876, N874, N239, N65, N156);
buf BUF1 (N877, N871);
nand NAND4 (N878, N849, N127, N657, N833);
and AND2 (N879, N877, N682);
xor XOR2 (N880, N876, N538);
nand NAND3 (N881, N870, N736, N445);
not NOT1 (N882, N872);
xor XOR2 (N883, N881, N85);
buf BUF1 (N884, N880);
not NOT1 (N885, N875);
and AND3 (N886, N878, N340, N535);
and AND4 (N887, N883, N402, N740, N704);
buf BUF1 (N888, N869);
buf BUF1 (N889, N882);
nand NAND3 (N890, N879, N531, N120);
buf BUF1 (N891, N845);
and AND2 (N892, N884, N618);
and AND4 (N893, N886, N235, N69, N447);
and AND2 (N894, N888, N136);
xor XOR2 (N895, N894, N655);
buf BUF1 (N896, N887);
nor NOR2 (N897, N896, N218);
not NOT1 (N898, N897);
and AND2 (N899, N895, N747);
or OR4 (N900, N891, N367, N97, N306);
nand NAND2 (N901, N898, N245);
not NOT1 (N902, N893);
nor NOR3 (N903, N890, N331, N347);
nand NAND3 (N904, N892, N422, N88);
xor XOR2 (N905, N904, N840);
xor XOR2 (N906, N835, N544);
nor NOR2 (N907, N885, N363);
nand NAND3 (N908, N902, N883, N52);
buf BUF1 (N909, N899);
and AND4 (N910, N908, N349, N42, N591);
nor NOR3 (N911, N903, N124, N726);
nor NOR3 (N912, N900, N373, N767);
and AND2 (N913, N910, N903);
nand NAND2 (N914, N913, N552);
nand NAND2 (N915, N901, N500);
or OR2 (N916, N915, N353);
and AND2 (N917, N889, N1);
nor NOR3 (N918, N868, N658, N532);
or OR3 (N919, N911, N498, N866);
nand NAND3 (N920, N905, N853, N113);
xor XOR2 (N921, N909, N319);
xor XOR2 (N922, N918, N424);
buf BUF1 (N923, N920);
buf BUF1 (N924, N923);
nand NAND2 (N925, N917, N635);
nand NAND2 (N926, N914, N506);
not NOT1 (N927, N907);
buf BUF1 (N928, N919);
and AND2 (N929, N916, N829);
xor XOR2 (N930, N925, N195);
and AND2 (N931, N922, N490);
buf BUF1 (N932, N927);
buf BUF1 (N933, N924);
not NOT1 (N934, N929);
not NOT1 (N935, N912);
or OR3 (N936, N935, N445, N555);
nand NAND2 (N937, N921, N171);
or OR2 (N938, N930, N893);
nand NAND4 (N939, N933, N784, N903, N625);
or OR2 (N940, N938, N258);
buf BUF1 (N941, N940);
buf BUF1 (N942, N936);
or OR2 (N943, N934, N844);
or OR4 (N944, N928, N34, N675, N398);
nor NOR4 (N945, N932, N809, N85, N113);
buf BUF1 (N946, N942);
not NOT1 (N947, N943);
nand NAND3 (N948, N941, N138, N504);
and AND2 (N949, N931, N478);
nor NOR3 (N950, N947, N841, N340);
buf BUF1 (N951, N945);
buf BUF1 (N952, N939);
buf BUF1 (N953, N950);
and AND4 (N954, N946, N339, N599, N611);
not NOT1 (N955, N953);
and AND3 (N956, N937, N507, N628);
xor XOR2 (N957, N951, N166);
or OR3 (N958, N954, N517, N282);
nor NOR4 (N959, N956, N509, N122, N450);
buf BUF1 (N960, N948);
xor XOR2 (N961, N944, N191);
and AND3 (N962, N926, N283, N607);
nand NAND2 (N963, N949, N509);
and AND4 (N964, N960, N511, N271, N41);
nor NOR3 (N965, N963, N393, N488);
nor NOR3 (N966, N952, N888, N235);
nand NAND2 (N967, N965, N59);
and AND3 (N968, N961, N179, N546);
nor NOR4 (N969, N959, N825, N424, N274);
nand NAND4 (N970, N964, N385, N328, N807);
buf BUF1 (N971, N966);
nor NOR4 (N972, N971, N327, N921, N76);
nand NAND2 (N973, N958, N882);
and AND2 (N974, N970, N62);
buf BUF1 (N975, N955);
and AND4 (N976, N962, N51, N850, N782);
and AND4 (N977, N968, N949, N133, N365);
and AND4 (N978, N973, N569, N778, N952);
xor XOR2 (N979, N976, N726);
and AND2 (N980, N972, N311);
nand NAND3 (N981, N957, N405, N729);
not NOT1 (N982, N969);
not NOT1 (N983, N978);
or OR4 (N984, N983, N342, N561, N58);
and AND2 (N985, N981, N91);
xor XOR2 (N986, N977, N864);
not NOT1 (N987, N906);
or OR3 (N988, N987, N40, N692);
buf BUF1 (N989, N975);
and AND4 (N990, N974, N907, N496, N213);
nor NOR2 (N991, N980, N440);
nor NOR4 (N992, N982, N985, N189, N647);
or OR3 (N993, N86, N390, N647);
xor XOR2 (N994, N990, N190);
buf BUF1 (N995, N994);
nand NAND2 (N996, N991, N537);
buf BUF1 (N997, N986);
not NOT1 (N998, N989);
nor NOR3 (N999, N995, N343, N312);
xor XOR2 (N1000, N993, N569);
xor XOR2 (N1001, N997, N110);
nor NOR2 (N1002, N998, N355);
nand NAND4 (N1003, N967, N426, N729, N337);
not NOT1 (N1004, N988);
nand NAND3 (N1005, N1000, N692, N242);
nor NOR3 (N1006, N1002, N931, N140);
and AND3 (N1007, N1003, N662, N631);
xor XOR2 (N1008, N984, N748);
not NOT1 (N1009, N999);
nor NOR2 (N1010, N992, N483);
and AND4 (N1011, N996, N533, N846, N560);
and AND2 (N1012, N1009, N782);
and AND3 (N1013, N1001, N30, N50);
or OR4 (N1014, N1012, N682, N123, N509);
nor NOR2 (N1015, N1004, N883);
not NOT1 (N1016, N1010);
not NOT1 (N1017, N1016);
xor XOR2 (N1018, N1007, N17);
not NOT1 (N1019, N1005);
nand NAND2 (N1020, N1011, N838);
nor NOR4 (N1021, N1017, N541, N646, N69);
nor NOR4 (N1022, N1013, N982, N376, N1019);
nand NAND2 (N1023, N358, N27);
not NOT1 (N1024, N979);
buf BUF1 (N1025, N1006);
xor XOR2 (N1026, N1025, N950);
buf BUF1 (N1027, N1020);
buf BUF1 (N1028, N1022);
or OR3 (N1029, N1028, N260, N902);
nand NAND2 (N1030, N1008, N273);
buf BUF1 (N1031, N1018);
or OR3 (N1032, N1023, N835, N538);
buf BUF1 (N1033, N1015);
buf BUF1 (N1034, N1024);
not NOT1 (N1035, N1031);
and AND4 (N1036, N1030, N224, N766, N491);
or OR3 (N1037, N1026, N862, N409);
not NOT1 (N1038, N1014);
nand NAND4 (N1039, N1033, N571, N607, N610);
and AND3 (N1040, N1036, N826, N998);
and AND3 (N1041, N1034, N327, N603);
not NOT1 (N1042, N1040);
and AND4 (N1043, N1039, N82, N136, N350);
nor NOR3 (N1044, N1037, N829, N685);
and AND3 (N1045, N1042, N843, N286);
or OR4 (N1046, N1041, N930, N812, N182);
buf BUF1 (N1047, N1035);
buf BUF1 (N1048, N1043);
and AND3 (N1049, N1038, N621, N911);
not NOT1 (N1050, N1048);
nor NOR4 (N1051, N1032, N747, N1027, N61);
and AND2 (N1052, N81, N381);
nand NAND2 (N1053, N1029, N320);
nand NAND2 (N1054, N1052, N633);
xor XOR2 (N1055, N1049, N380);
not NOT1 (N1056, N1053);
buf BUF1 (N1057, N1055);
xor XOR2 (N1058, N1057, N95);
xor XOR2 (N1059, N1058, N701);
not NOT1 (N1060, N1056);
nand NAND2 (N1061, N1059, N296);
nand NAND2 (N1062, N1045, N123);
buf BUF1 (N1063, N1051);
not NOT1 (N1064, N1050);
and AND4 (N1065, N1064, N656, N256, N246);
not NOT1 (N1066, N1044);
nor NOR2 (N1067, N1062, N222);
nor NOR3 (N1068, N1021, N183, N297);
xor XOR2 (N1069, N1067, N573);
buf BUF1 (N1070, N1066);
and AND4 (N1071, N1060, N687, N368, N769);
and AND3 (N1072, N1063, N275, N673);
buf BUF1 (N1073, N1071);
and AND2 (N1074, N1061, N806);
nand NAND3 (N1075, N1068, N162, N492);
nand NAND4 (N1076, N1054, N841, N681, N788);
and AND2 (N1077, N1047, N543);
buf BUF1 (N1078, N1072);
nor NOR2 (N1079, N1070, N102);
or OR2 (N1080, N1065, N358);
nand NAND3 (N1081, N1074, N135, N406);
nor NOR3 (N1082, N1046, N170, N885);
xor XOR2 (N1083, N1076, N180);
and AND2 (N1084, N1075, N338);
nand NAND3 (N1085, N1079, N994, N488);
nor NOR2 (N1086, N1084, N951);
and AND2 (N1087, N1078, N594);
xor XOR2 (N1088, N1083, N691);
xor XOR2 (N1089, N1085, N716);
not NOT1 (N1090, N1088);
not NOT1 (N1091, N1087);
nand NAND3 (N1092, N1090, N1007, N776);
nor NOR3 (N1093, N1089, N400, N916);
not NOT1 (N1094, N1077);
xor XOR2 (N1095, N1091, N650);
not NOT1 (N1096, N1081);
and AND2 (N1097, N1086, N48);
not NOT1 (N1098, N1097);
and AND2 (N1099, N1080, N56);
buf BUF1 (N1100, N1082);
buf BUF1 (N1101, N1099);
nand NAND4 (N1102, N1069, N320, N159, N545);
and AND3 (N1103, N1093, N138, N503);
buf BUF1 (N1104, N1100);
xor XOR2 (N1105, N1103, N404);
buf BUF1 (N1106, N1098);
nand NAND2 (N1107, N1101, N491);
xor XOR2 (N1108, N1096, N366);
or OR4 (N1109, N1094, N42, N709, N761);
not NOT1 (N1110, N1104);
buf BUF1 (N1111, N1109);
buf BUF1 (N1112, N1111);
not NOT1 (N1113, N1095);
nand NAND3 (N1114, N1092, N1015, N548);
nor NOR2 (N1115, N1113, N688);
nor NOR2 (N1116, N1102, N1086);
and AND2 (N1117, N1114, N851);
nand NAND4 (N1118, N1073, N1116, N582, N366);
or OR2 (N1119, N391, N455);
nand NAND4 (N1120, N1119, N789, N769, N917);
xor XOR2 (N1121, N1117, N482);
nor NOR4 (N1122, N1112, N490, N767, N927);
nor NOR4 (N1123, N1120, N640, N1108, N404);
not NOT1 (N1124, N1057);
nand NAND3 (N1125, N1106, N48, N1040);
nor NOR3 (N1126, N1105, N111, N975);
nand NAND3 (N1127, N1107, N228, N85);
and AND3 (N1128, N1122, N953, N543);
nor NOR2 (N1129, N1126, N515);
nand NAND3 (N1130, N1129, N427, N405);
buf BUF1 (N1131, N1124);
nor NOR2 (N1132, N1125, N147);
buf BUF1 (N1133, N1121);
and AND3 (N1134, N1110, N545, N997);
or OR4 (N1135, N1130, N983, N977, N119);
not NOT1 (N1136, N1127);
nor NOR2 (N1137, N1136, N238);
nor NOR3 (N1138, N1132, N191, N395);
nor NOR3 (N1139, N1118, N766, N271);
not NOT1 (N1140, N1138);
buf BUF1 (N1141, N1123);
nand NAND2 (N1142, N1139, N281);
not NOT1 (N1143, N1142);
or OR3 (N1144, N1128, N934, N887);
xor XOR2 (N1145, N1135, N341);
xor XOR2 (N1146, N1115, N113);
not NOT1 (N1147, N1140);
nor NOR4 (N1148, N1137, N190, N684, N8);
xor XOR2 (N1149, N1144, N641);
not NOT1 (N1150, N1143);
or OR4 (N1151, N1141, N365, N792, N860);
not NOT1 (N1152, N1146);
or OR4 (N1153, N1150, N901, N187, N680);
nand NAND3 (N1154, N1131, N958, N344);
and AND3 (N1155, N1134, N1153, N914);
and AND3 (N1156, N320, N287, N814);
xor XOR2 (N1157, N1155, N325);
nor NOR3 (N1158, N1145, N792, N322);
nand NAND3 (N1159, N1148, N464, N272);
xor XOR2 (N1160, N1133, N153);
buf BUF1 (N1161, N1156);
buf BUF1 (N1162, N1152);
or OR2 (N1163, N1158, N843);
and AND2 (N1164, N1157, N617);
nand NAND3 (N1165, N1163, N201, N985);
nor NOR4 (N1166, N1161, N439, N1004, N85);
xor XOR2 (N1167, N1162, N306);
buf BUF1 (N1168, N1149);
or OR3 (N1169, N1168, N930, N58);
xor XOR2 (N1170, N1154, N1138);
nor NOR4 (N1171, N1167, N1084, N726, N366);
or OR3 (N1172, N1170, N505, N155);
and AND4 (N1173, N1147, N30, N931, N1137);
nand NAND3 (N1174, N1171, N225, N106);
buf BUF1 (N1175, N1165);
nand NAND4 (N1176, N1174, N727, N618, N695);
not NOT1 (N1177, N1160);
not NOT1 (N1178, N1176);
not NOT1 (N1179, N1178);
nor NOR2 (N1180, N1166, N281);
or OR2 (N1181, N1179, N808);
xor XOR2 (N1182, N1180, N890);
or OR2 (N1183, N1181, N478);
nor NOR2 (N1184, N1177, N464);
and AND3 (N1185, N1184, N240, N819);
nand NAND3 (N1186, N1175, N404, N326);
not NOT1 (N1187, N1169);
xor XOR2 (N1188, N1183, N917);
and AND3 (N1189, N1173, N3, N742);
or OR4 (N1190, N1186, N278, N1096, N144);
or OR4 (N1191, N1190, N1167, N122, N127);
xor XOR2 (N1192, N1164, N545);
nand NAND4 (N1193, N1191, N746, N1017, N1180);
or OR3 (N1194, N1185, N71, N175);
not NOT1 (N1195, N1189);
xor XOR2 (N1196, N1192, N30);
xor XOR2 (N1197, N1188, N908);
xor XOR2 (N1198, N1194, N1180);
or OR2 (N1199, N1159, N354);
xor XOR2 (N1200, N1151, N417);
nor NOR2 (N1201, N1198, N459);
buf BUF1 (N1202, N1187);
not NOT1 (N1203, N1193);
nand NAND3 (N1204, N1203, N820, N300);
buf BUF1 (N1205, N1204);
xor XOR2 (N1206, N1201, N585);
buf BUF1 (N1207, N1205);
and AND3 (N1208, N1172, N456, N110);
buf BUF1 (N1209, N1207);
not NOT1 (N1210, N1208);
buf BUF1 (N1211, N1210);
xor XOR2 (N1212, N1199, N1205);
not NOT1 (N1213, N1200);
or OR2 (N1214, N1213, N32);
and AND2 (N1215, N1206, N400);
nor NOR3 (N1216, N1182, N131, N36);
or OR2 (N1217, N1202, N497);
or OR2 (N1218, N1211, N1171);
nor NOR3 (N1219, N1215, N822, N679);
nand NAND2 (N1220, N1195, N1153);
buf BUF1 (N1221, N1209);
xor XOR2 (N1222, N1216, N256);
buf BUF1 (N1223, N1217);
and AND2 (N1224, N1221, N457);
buf BUF1 (N1225, N1196);
nand NAND2 (N1226, N1214, N363);
and AND2 (N1227, N1218, N135);
and AND3 (N1228, N1224, N100, N288);
xor XOR2 (N1229, N1225, N494);
and AND3 (N1230, N1229, N361, N443);
not NOT1 (N1231, N1228);
or OR2 (N1232, N1197, N495);
nor NOR3 (N1233, N1220, N376, N399);
xor XOR2 (N1234, N1232, N701);
not NOT1 (N1235, N1230);
and AND3 (N1236, N1234, N501, N1018);
nand NAND3 (N1237, N1226, N76, N48);
xor XOR2 (N1238, N1212, N700);
or OR2 (N1239, N1219, N383);
and AND2 (N1240, N1231, N353);
xor XOR2 (N1241, N1239, N670);
buf BUF1 (N1242, N1223);
xor XOR2 (N1243, N1237, N753);
buf BUF1 (N1244, N1233);
or OR4 (N1245, N1235, N893, N700, N16);
and AND2 (N1246, N1238, N388);
xor XOR2 (N1247, N1244, N357);
xor XOR2 (N1248, N1241, N35);
nand NAND3 (N1249, N1240, N1116, N812);
nand NAND3 (N1250, N1227, N174, N56);
not NOT1 (N1251, N1249);
and AND3 (N1252, N1242, N711, N623);
and AND3 (N1253, N1243, N1209, N1187);
xor XOR2 (N1254, N1245, N428);
and AND2 (N1255, N1247, N1090);
nand NAND2 (N1256, N1252, N624);
or OR3 (N1257, N1251, N922, N1177);
buf BUF1 (N1258, N1254);
nand NAND4 (N1259, N1236, N811, N95, N950);
nor NOR4 (N1260, N1259, N750, N851, N1165);
and AND4 (N1261, N1246, N735, N1114, N33);
xor XOR2 (N1262, N1248, N1050);
and AND4 (N1263, N1261, N378, N751, N1164);
buf BUF1 (N1264, N1250);
xor XOR2 (N1265, N1257, N233);
nand NAND4 (N1266, N1264, N644, N404, N1197);
or OR2 (N1267, N1255, N165);
and AND4 (N1268, N1222, N757, N1032, N614);
not NOT1 (N1269, N1253);
nor NOR3 (N1270, N1269, N366, N939);
nand NAND4 (N1271, N1268, N92, N371, N520);
or OR2 (N1272, N1260, N710);
and AND2 (N1273, N1258, N672);
or OR2 (N1274, N1256, N126);
nor NOR3 (N1275, N1265, N912, N534);
nor NOR3 (N1276, N1267, N270, N240);
buf BUF1 (N1277, N1275);
not NOT1 (N1278, N1274);
xor XOR2 (N1279, N1262, N738);
xor XOR2 (N1280, N1271, N258);
and AND4 (N1281, N1276, N1234, N419, N147);
buf BUF1 (N1282, N1270);
not NOT1 (N1283, N1282);
nor NOR4 (N1284, N1266, N331, N854, N1068);
buf BUF1 (N1285, N1263);
xor XOR2 (N1286, N1279, N683);
nand NAND4 (N1287, N1277, N228, N1066, N742);
nor NOR2 (N1288, N1287, N557);
and AND3 (N1289, N1278, N506, N189);
not NOT1 (N1290, N1281);
nand NAND2 (N1291, N1284, N15);
xor XOR2 (N1292, N1290, N878);
nand NAND3 (N1293, N1273, N210, N271);
or OR2 (N1294, N1291, N244);
and AND4 (N1295, N1272, N589, N770, N858);
not NOT1 (N1296, N1288);
xor XOR2 (N1297, N1293, N685);
or OR3 (N1298, N1285, N721, N1037);
nand NAND3 (N1299, N1280, N388, N153);
nor NOR3 (N1300, N1295, N795, N1253);
nor NOR3 (N1301, N1286, N198, N332);
buf BUF1 (N1302, N1296);
nor NOR3 (N1303, N1302, N110, N97);
nand NAND3 (N1304, N1289, N1153, N496);
or OR2 (N1305, N1297, N1040);
not NOT1 (N1306, N1292);
xor XOR2 (N1307, N1294, N413);
buf BUF1 (N1308, N1299);
nor NOR4 (N1309, N1303, N1308, N286, N628);
nand NAND4 (N1310, N526, N1186, N394, N398);
not NOT1 (N1311, N1310);
buf BUF1 (N1312, N1301);
xor XOR2 (N1313, N1311, N498);
not NOT1 (N1314, N1306);
xor XOR2 (N1315, N1305, N767);
xor XOR2 (N1316, N1312, N1222);
and AND4 (N1317, N1313, N161, N587, N679);
not NOT1 (N1318, N1300);
buf BUF1 (N1319, N1298);
not NOT1 (N1320, N1316);
or OR3 (N1321, N1317, N204, N490);
not NOT1 (N1322, N1315);
xor XOR2 (N1323, N1307, N435);
xor XOR2 (N1324, N1320, N346);
nand NAND3 (N1325, N1304, N1059, N220);
nand NAND3 (N1326, N1314, N649, N935);
buf BUF1 (N1327, N1325);
nand NAND2 (N1328, N1319, N1009);
nor NOR4 (N1329, N1283, N890, N128, N708);
xor XOR2 (N1330, N1324, N798);
nand NAND3 (N1331, N1321, N393, N287);
not NOT1 (N1332, N1318);
buf BUF1 (N1333, N1329);
nor NOR2 (N1334, N1323, N476);
xor XOR2 (N1335, N1322, N491);
and AND3 (N1336, N1330, N886, N319);
and AND3 (N1337, N1333, N109, N1052);
nor NOR4 (N1338, N1327, N629, N680, N78);
and AND2 (N1339, N1332, N898);
nand NAND3 (N1340, N1339, N519, N56);
and AND3 (N1341, N1336, N262, N743);
or OR4 (N1342, N1334, N162, N493, N159);
not NOT1 (N1343, N1338);
not NOT1 (N1344, N1343);
buf BUF1 (N1345, N1335);
nor NOR3 (N1346, N1344, N420, N1272);
nand NAND2 (N1347, N1342, N856);
nor NOR2 (N1348, N1328, N1206);
or OR2 (N1349, N1348, N1172);
xor XOR2 (N1350, N1340, N1337);
xor XOR2 (N1351, N604, N175);
not NOT1 (N1352, N1350);
or OR4 (N1353, N1352, N476, N547, N294);
nor NOR4 (N1354, N1341, N117, N1341, N47);
xor XOR2 (N1355, N1346, N491);
nor NOR2 (N1356, N1355, N1345);
or OR4 (N1357, N225, N773, N1092, N448);
nor NOR2 (N1358, N1309, N514);
not NOT1 (N1359, N1358);
not NOT1 (N1360, N1326);
not NOT1 (N1361, N1360);
buf BUF1 (N1362, N1349);
buf BUF1 (N1363, N1331);
or OR4 (N1364, N1357, N721, N593, N940);
or OR2 (N1365, N1356, N1029);
nor NOR4 (N1366, N1347, N558, N87, N431);
nand NAND2 (N1367, N1366, N342);
xor XOR2 (N1368, N1353, N551);
or OR2 (N1369, N1362, N411);
not NOT1 (N1370, N1367);
nand NAND4 (N1371, N1364, N259, N1243, N177);
nand NAND2 (N1372, N1359, N184);
nand NAND4 (N1373, N1369, N315, N1177, N1089);
or OR3 (N1374, N1371, N1188, N1135);
or OR3 (N1375, N1374, N1101, N740);
and AND4 (N1376, N1368, N927, N361, N236);
xor XOR2 (N1377, N1376, N1180);
xor XOR2 (N1378, N1377, N816);
nand NAND3 (N1379, N1365, N808, N260);
nor NOR3 (N1380, N1373, N414, N1352);
nor NOR4 (N1381, N1378, N1076, N994, N359);
nand NAND3 (N1382, N1361, N73, N13);
nand NAND2 (N1383, N1351, N1005);
not NOT1 (N1384, N1379);
nand NAND4 (N1385, N1382, N1192, N1146, N944);
not NOT1 (N1386, N1363);
not NOT1 (N1387, N1385);
and AND2 (N1388, N1387, N332);
nand NAND2 (N1389, N1388, N426);
and AND3 (N1390, N1375, N1021, N729);
and AND4 (N1391, N1386, N500, N106, N1192);
and AND4 (N1392, N1391, N707, N813, N337);
xor XOR2 (N1393, N1384, N192);
xor XOR2 (N1394, N1393, N1061);
or OR4 (N1395, N1381, N910, N1271, N991);
not NOT1 (N1396, N1380);
xor XOR2 (N1397, N1395, N812);
nor NOR3 (N1398, N1354, N444, N178);
buf BUF1 (N1399, N1394);
not NOT1 (N1400, N1392);
nor NOR3 (N1401, N1400, N222, N172);
or OR2 (N1402, N1389, N465);
xor XOR2 (N1403, N1398, N966);
and AND4 (N1404, N1372, N102, N1226, N554);
buf BUF1 (N1405, N1397);
buf BUF1 (N1406, N1404);
xor XOR2 (N1407, N1370, N193);
xor XOR2 (N1408, N1390, N427);
or OR3 (N1409, N1396, N682, N218);
nand NAND3 (N1410, N1383, N360, N262);
nor NOR3 (N1411, N1402, N981, N789);
and AND3 (N1412, N1411, N1367, N994);
xor XOR2 (N1413, N1399, N174);
or OR2 (N1414, N1410, N1249);
buf BUF1 (N1415, N1412);
xor XOR2 (N1416, N1405, N1180);
nor NOR4 (N1417, N1406, N565, N548, N1328);
nor NOR4 (N1418, N1416, N66, N1373, N585);
xor XOR2 (N1419, N1417, N486);
nor NOR3 (N1420, N1401, N28, N624);
buf BUF1 (N1421, N1403);
not NOT1 (N1422, N1418);
or OR3 (N1423, N1407, N1209, N1012);
nor NOR2 (N1424, N1408, N153);
buf BUF1 (N1425, N1414);
nor NOR2 (N1426, N1424, N752);
nand NAND2 (N1427, N1415, N683);
not NOT1 (N1428, N1422);
and AND2 (N1429, N1423, N1102);
nor NOR3 (N1430, N1427, N243, N112);
not NOT1 (N1431, N1425);
nand NAND3 (N1432, N1426, N1145, N130);
and AND2 (N1433, N1431, N486);
buf BUF1 (N1434, N1432);
and AND4 (N1435, N1433, N454, N1219, N64);
or OR3 (N1436, N1409, N817, N1345);
xor XOR2 (N1437, N1421, N233);
and AND2 (N1438, N1419, N355);
buf BUF1 (N1439, N1434);
nor NOR3 (N1440, N1429, N1008, N318);
nor NOR4 (N1441, N1430, N713, N1350, N473);
or OR3 (N1442, N1438, N1175, N1334);
nor NOR2 (N1443, N1413, N894);
xor XOR2 (N1444, N1439, N231);
nor NOR3 (N1445, N1440, N17, N429);
nand NAND2 (N1446, N1420, N909);
nand NAND2 (N1447, N1442, N520);
and AND4 (N1448, N1445, N1222, N523, N1071);
nor NOR2 (N1449, N1446, N783);
nor NOR4 (N1450, N1444, N536, N561, N546);
buf BUF1 (N1451, N1448);
buf BUF1 (N1452, N1428);
not NOT1 (N1453, N1443);
buf BUF1 (N1454, N1450);
buf BUF1 (N1455, N1435);
nand NAND3 (N1456, N1452, N778, N153);
nand NAND4 (N1457, N1447, N1346, N422, N327);
buf BUF1 (N1458, N1449);
not NOT1 (N1459, N1436);
not NOT1 (N1460, N1441);
xor XOR2 (N1461, N1453, N1111);
not NOT1 (N1462, N1459);
not NOT1 (N1463, N1458);
xor XOR2 (N1464, N1451, N378);
buf BUF1 (N1465, N1457);
nor NOR2 (N1466, N1463, N941);
buf BUF1 (N1467, N1460);
or OR2 (N1468, N1462, N12);
not NOT1 (N1469, N1454);
and AND4 (N1470, N1456, N392, N802, N948);
nand NAND2 (N1471, N1461, N269);
nor NOR3 (N1472, N1466, N23, N1435);
nor NOR4 (N1473, N1437, N847, N118, N544);
buf BUF1 (N1474, N1470);
buf BUF1 (N1475, N1455);
xor XOR2 (N1476, N1469, N1143);
nor NOR4 (N1477, N1475, N676, N1424, N317);
nand NAND2 (N1478, N1476, N684);
or OR4 (N1479, N1468, N105, N621, N125);
nor NOR2 (N1480, N1465, N1120);
nor NOR4 (N1481, N1480, N656, N1086, N18);
nor NOR3 (N1482, N1472, N560, N1395);
not NOT1 (N1483, N1477);
and AND3 (N1484, N1473, N1469, N617);
buf BUF1 (N1485, N1481);
nor NOR2 (N1486, N1479, N88);
buf BUF1 (N1487, N1483);
or OR4 (N1488, N1486, N1180, N234, N283);
or OR4 (N1489, N1482, N1326, N944, N402);
or OR2 (N1490, N1464, N255);
not NOT1 (N1491, N1489);
not NOT1 (N1492, N1491);
nand NAND2 (N1493, N1471, N1205);
nand NAND3 (N1494, N1478, N225, N1095);
not NOT1 (N1495, N1467);
nor NOR3 (N1496, N1494, N50, N562);
or OR4 (N1497, N1487, N775, N1173, N587);
nand NAND2 (N1498, N1497, N1094);
or OR2 (N1499, N1488, N28);
not NOT1 (N1500, N1485);
buf BUF1 (N1501, N1474);
or OR2 (N1502, N1490, N1311);
not NOT1 (N1503, N1492);
and AND2 (N1504, N1496, N781);
not NOT1 (N1505, N1501);
nand NAND4 (N1506, N1484, N736, N1336, N907);
nand NAND3 (N1507, N1498, N514, N613);
nor NOR3 (N1508, N1504, N1425, N789);
or OR4 (N1509, N1495, N398, N1357, N584);
nor NOR3 (N1510, N1493, N586, N202);
or OR4 (N1511, N1503, N729, N370, N837);
or OR4 (N1512, N1505, N1231, N1099, N1473);
nor NOR4 (N1513, N1499, N315, N1158, N173);
buf BUF1 (N1514, N1512);
nand NAND4 (N1515, N1506, N1064, N537, N1377);
not NOT1 (N1516, N1507);
xor XOR2 (N1517, N1511, N1413);
not NOT1 (N1518, N1517);
not NOT1 (N1519, N1510);
not NOT1 (N1520, N1518);
or OR3 (N1521, N1502, N1128, N873);
nand NAND2 (N1522, N1508, N1439);
buf BUF1 (N1523, N1515);
or OR2 (N1524, N1519, N590);
or OR3 (N1525, N1513, N1149, N1163);
nand NAND3 (N1526, N1520, N1205, N300);
or OR2 (N1527, N1516, N666);
nand NAND4 (N1528, N1527, N1007, N173, N304);
xor XOR2 (N1529, N1526, N589);
or OR4 (N1530, N1523, N1402, N180, N854);
not NOT1 (N1531, N1525);
or OR3 (N1532, N1528, N281, N1520);
and AND4 (N1533, N1509, N710, N780, N1424);
not NOT1 (N1534, N1532);
nor NOR2 (N1535, N1531, N895);
or OR3 (N1536, N1530, N257, N1468);
or OR2 (N1537, N1534, N1313);
nand NAND4 (N1538, N1529, N526, N1295, N259);
nand NAND3 (N1539, N1521, N439, N649);
xor XOR2 (N1540, N1524, N1174);
and AND4 (N1541, N1533, N945, N1111, N154);
or OR2 (N1542, N1514, N129);
nand NAND3 (N1543, N1542, N1008, N1143);
buf BUF1 (N1544, N1500);
buf BUF1 (N1545, N1538);
nor NOR4 (N1546, N1541, N429, N1030, N186);
xor XOR2 (N1547, N1545, N1076);
and AND2 (N1548, N1536, N860);
not NOT1 (N1549, N1543);
not NOT1 (N1550, N1549);
nand NAND3 (N1551, N1546, N1379, N736);
buf BUF1 (N1552, N1540);
or OR3 (N1553, N1551, N300, N965);
buf BUF1 (N1554, N1548);
or OR4 (N1555, N1544, N84, N211, N1498);
buf BUF1 (N1556, N1554);
nor NOR3 (N1557, N1535, N285, N1233);
nor NOR2 (N1558, N1547, N1268);
or OR3 (N1559, N1556, N1534, N1392);
not NOT1 (N1560, N1558);
not NOT1 (N1561, N1559);
xor XOR2 (N1562, N1560, N1475);
nor NOR3 (N1563, N1555, N730, N651);
xor XOR2 (N1564, N1522, N630);
nand NAND2 (N1565, N1564, N911);
nor NOR3 (N1566, N1557, N1031, N75);
nand NAND2 (N1567, N1561, N531);
or OR2 (N1568, N1562, N482);
and AND3 (N1569, N1567, N692, N1014);
xor XOR2 (N1570, N1553, N51);
or OR3 (N1571, N1563, N690, N363);
nor NOR3 (N1572, N1537, N307, N488);
buf BUF1 (N1573, N1572);
nand NAND2 (N1574, N1565, N1317);
nand NAND3 (N1575, N1550, N1565, N1016);
buf BUF1 (N1576, N1568);
nor NOR4 (N1577, N1566, N166, N447, N470);
xor XOR2 (N1578, N1577, N1377);
and AND2 (N1579, N1570, N334);
xor XOR2 (N1580, N1574, N303);
buf BUF1 (N1581, N1571);
nor NOR4 (N1582, N1552, N19, N1186, N656);
nor NOR3 (N1583, N1580, N1483, N102);
nand NAND3 (N1584, N1578, N205, N366);
nand NAND3 (N1585, N1584, N869, N698);
nand NAND4 (N1586, N1579, N835, N1455, N1193);
nand NAND2 (N1587, N1539, N1422);
or OR3 (N1588, N1581, N720, N1243);
buf BUF1 (N1589, N1586);
buf BUF1 (N1590, N1569);
xor XOR2 (N1591, N1575, N850);
xor XOR2 (N1592, N1591, N990);
and AND4 (N1593, N1588, N1349, N1589, N1162);
nor NOR2 (N1594, N1447, N239);
xor XOR2 (N1595, N1585, N262);
xor XOR2 (N1596, N1594, N621);
and AND2 (N1597, N1587, N1191);
nand NAND3 (N1598, N1592, N414, N1095);
buf BUF1 (N1599, N1596);
or OR2 (N1600, N1598, N26);
buf BUF1 (N1601, N1595);
xor XOR2 (N1602, N1597, N540);
nand NAND4 (N1603, N1593, N14, N374, N132);
xor XOR2 (N1604, N1599, N971);
or OR2 (N1605, N1573, N663);
or OR2 (N1606, N1601, N351);
not NOT1 (N1607, N1602);
nor NOR3 (N1608, N1605, N540, N39);
nor NOR2 (N1609, N1576, N1222);
not NOT1 (N1610, N1603);
not NOT1 (N1611, N1606);
not NOT1 (N1612, N1607);
or OR2 (N1613, N1582, N103);
or OR2 (N1614, N1610, N690);
buf BUF1 (N1615, N1600);
and AND3 (N1616, N1615, N1500, N742);
not NOT1 (N1617, N1590);
and AND3 (N1618, N1604, N458, N335);
nand NAND4 (N1619, N1611, N704, N233, N1436);
or OR4 (N1620, N1616, N1080, N669, N241);
not NOT1 (N1621, N1620);
or OR2 (N1622, N1619, N497);
nor NOR4 (N1623, N1612, N1106, N1539, N347);
xor XOR2 (N1624, N1583, N1044);
not NOT1 (N1625, N1624);
nor NOR3 (N1626, N1625, N1396, N600);
nand NAND3 (N1627, N1609, N744, N616);
or OR3 (N1628, N1608, N1229, N240);
nand NAND2 (N1629, N1613, N455);
or OR4 (N1630, N1614, N698, N177, N166);
xor XOR2 (N1631, N1629, N1605);
nand NAND2 (N1632, N1621, N1091);
nor NOR4 (N1633, N1618, N1209, N1600, N1091);
nand NAND3 (N1634, N1630, N734, N774);
nor NOR4 (N1635, N1626, N494, N1043, N1512);
or OR2 (N1636, N1633, N492);
or OR3 (N1637, N1617, N1198, N789);
and AND4 (N1638, N1636, N1511, N422, N1398);
and AND2 (N1639, N1623, N446);
buf BUF1 (N1640, N1622);
or OR4 (N1641, N1639, N34, N836, N748);
nor NOR3 (N1642, N1641, N1251, N1332);
or OR2 (N1643, N1642, N596);
buf BUF1 (N1644, N1631);
or OR3 (N1645, N1634, N90, N719);
or OR3 (N1646, N1640, N771, N224);
xor XOR2 (N1647, N1635, N162);
buf BUF1 (N1648, N1638);
nand NAND2 (N1649, N1644, N1269);
nand NAND4 (N1650, N1632, N1170, N1213, N261);
not NOT1 (N1651, N1650);
buf BUF1 (N1652, N1628);
buf BUF1 (N1653, N1647);
or OR2 (N1654, N1637, N1096);
xor XOR2 (N1655, N1649, N642);
nand NAND4 (N1656, N1653, N391, N1339, N747);
xor XOR2 (N1657, N1646, N805);
xor XOR2 (N1658, N1643, N465);
nand NAND3 (N1659, N1652, N14, N1520);
xor XOR2 (N1660, N1645, N622);
xor XOR2 (N1661, N1656, N1500);
or OR3 (N1662, N1655, N1263, N1472);
nor NOR4 (N1663, N1651, N358, N1557, N502);
buf BUF1 (N1664, N1662);
nand NAND2 (N1665, N1664, N1021);
xor XOR2 (N1666, N1659, N1185);
or OR2 (N1667, N1661, N1215);
nand NAND2 (N1668, N1658, N1162);
nor NOR3 (N1669, N1654, N25, N1315);
nand NAND4 (N1670, N1648, N584, N293, N732);
nand NAND3 (N1671, N1666, N382, N367);
not NOT1 (N1672, N1669);
xor XOR2 (N1673, N1660, N783);
or OR2 (N1674, N1627, N1627);
and AND2 (N1675, N1671, N606);
xor XOR2 (N1676, N1674, N803);
nor NOR4 (N1677, N1665, N820, N1048, N600);
nand NAND2 (N1678, N1657, N360);
not NOT1 (N1679, N1673);
buf BUF1 (N1680, N1676);
or OR4 (N1681, N1678, N502, N1002, N173);
buf BUF1 (N1682, N1679);
not NOT1 (N1683, N1668);
buf BUF1 (N1684, N1681);
and AND2 (N1685, N1663, N849);
nor NOR2 (N1686, N1684, N1214);
not NOT1 (N1687, N1677);
or OR3 (N1688, N1687, N344, N814);
xor XOR2 (N1689, N1683, N667);
not NOT1 (N1690, N1689);
xor XOR2 (N1691, N1686, N1148);
not NOT1 (N1692, N1670);
nor NOR3 (N1693, N1685, N299, N981);
nor NOR4 (N1694, N1693, N778, N463, N1037);
buf BUF1 (N1695, N1694);
or OR3 (N1696, N1691, N1493, N891);
xor XOR2 (N1697, N1672, N573);
nand NAND3 (N1698, N1692, N1037, N436);
xor XOR2 (N1699, N1698, N350);
buf BUF1 (N1700, N1696);
nor NOR2 (N1701, N1682, N1478);
xor XOR2 (N1702, N1688, N1485);
nand NAND4 (N1703, N1699, N1321, N354, N902);
or OR4 (N1704, N1702, N688, N1045, N532);
xor XOR2 (N1705, N1680, N860);
buf BUF1 (N1706, N1704);
nand NAND4 (N1707, N1675, N1312, N1244, N588);
buf BUF1 (N1708, N1697);
xor XOR2 (N1709, N1706, N587);
and AND2 (N1710, N1703, N756);
xor XOR2 (N1711, N1700, N228);
nand NAND3 (N1712, N1705, N836, N876);
and AND2 (N1713, N1667, N378);
buf BUF1 (N1714, N1708);
or OR2 (N1715, N1709, N1547);
and AND3 (N1716, N1714, N1298, N206);
nor NOR2 (N1717, N1716, N274);
not NOT1 (N1718, N1713);
not NOT1 (N1719, N1695);
nor NOR3 (N1720, N1715, N468, N655);
nand NAND2 (N1721, N1717, N1164);
nand NAND2 (N1722, N1712, N1245);
nand NAND3 (N1723, N1711, N236, N1562);
xor XOR2 (N1724, N1701, N208);
not NOT1 (N1725, N1719);
buf BUF1 (N1726, N1720);
not NOT1 (N1727, N1722);
and AND3 (N1728, N1710, N1029, N1049);
nor NOR3 (N1729, N1727, N1309, N785);
or OR2 (N1730, N1721, N863);
and AND2 (N1731, N1690, N434);
and AND4 (N1732, N1730, N1454, N590, N1707);
or OR4 (N1733, N500, N975, N602, N528);
nand NAND3 (N1734, N1733, N1008, N819);
or OR4 (N1735, N1725, N304, N187, N1440);
buf BUF1 (N1736, N1734);
nor NOR4 (N1737, N1718, N529, N745, N1475);
xor XOR2 (N1738, N1732, N1068);
and AND2 (N1739, N1737, N1690);
buf BUF1 (N1740, N1736);
nor NOR3 (N1741, N1724, N747, N1605);
nand NAND2 (N1742, N1740, N963);
not NOT1 (N1743, N1738);
not NOT1 (N1744, N1729);
nand NAND2 (N1745, N1739, N895);
nand NAND4 (N1746, N1723, N212, N1226, N1604);
nand NAND2 (N1747, N1743, N972);
not NOT1 (N1748, N1728);
nor NOR2 (N1749, N1741, N1660);
nand NAND2 (N1750, N1744, N1391);
or OR4 (N1751, N1735, N986, N644, N824);
buf BUF1 (N1752, N1731);
and AND3 (N1753, N1750, N159, N218);
and AND3 (N1754, N1726, N747, N1415);
nand NAND3 (N1755, N1752, N206, N1152);
xor XOR2 (N1756, N1742, N1698);
not NOT1 (N1757, N1753);
buf BUF1 (N1758, N1745);
or OR2 (N1759, N1754, N50);
not NOT1 (N1760, N1759);
buf BUF1 (N1761, N1749);
not NOT1 (N1762, N1746);
xor XOR2 (N1763, N1757, N417);
xor XOR2 (N1764, N1756, N660);
or OR3 (N1765, N1755, N1752, N982);
and AND4 (N1766, N1762, N1386, N1541, N657);
nand NAND3 (N1767, N1751, N853, N376);
xor XOR2 (N1768, N1747, N728);
buf BUF1 (N1769, N1764);
not NOT1 (N1770, N1761);
buf BUF1 (N1771, N1758);
xor XOR2 (N1772, N1769, N1007);
nor NOR2 (N1773, N1760, N1431);
or OR4 (N1774, N1763, N869, N1508, N312);
xor XOR2 (N1775, N1772, N502);
xor XOR2 (N1776, N1770, N707);
nand NAND3 (N1777, N1776, N56, N610);
nand NAND2 (N1778, N1777, N1259);
nand NAND4 (N1779, N1768, N1553, N703, N72);
nand NAND3 (N1780, N1774, N1335, N498);
nor NOR4 (N1781, N1780, N78, N131, N795);
buf BUF1 (N1782, N1778);
buf BUF1 (N1783, N1782);
or OR3 (N1784, N1773, N771, N849);
nor NOR2 (N1785, N1767, N211);
buf BUF1 (N1786, N1781);
and AND2 (N1787, N1775, N50);
or OR2 (N1788, N1784, N1460);
xor XOR2 (N1789, N1748, N766);
nand NAND4 (N1790, N1786, N898, N1753, N127);
or OR3 (N1791, N1771, N263, N1120);
and AND4 (N1792, N1765, N323, N1076, N1340);
not NOT1 (N1793, N1787);
nor NOR2 (N1794, N1793, N1219);
buf BUF1 (N1795, N1792);
nor NOR4 (N1796, N1790, N19, N380, N1671);
not NOT1 (N1797, N1789);
buf BUF1 (N1798, N1797);
and AND4 (N1799, N1785, N232, N523, N366);
and AND2 (N1800, N1794, N489);
and AND4 (N1801, N1798, N757, N1695, N10);
nand NAND3 (N1802, N1796, N1657, N575);
not NOT1 (N1803, N1801);
buf BUF1 (N1804, N1783);
xor XOR2 (N1805, N1766, N1620);
xor XOR2 (N1806, N1791, N1717);
nand NAND4 (N1807, N1800, N1203, N1165, N1495);
nand NAND4 (N1808, N1806, N1466, N1269, N1684);
xor XOR2 (N1809, N1788, N253);
xor XOR2 (N1810, N1799, N420);
buf BUF1 (N1811, N1810);
or OR4 (N1812, N1811, N1790, N125, N1742);
nor NOR4 (N1813, N1809, N439, N1696, N236);
or OR4 (N1814, N1804, N498, N519, N1302);
nor NOR2 (N1815, N1808, N1694);
buf BUF1 (N1816, N1805);
or OR3 (N1817, N1802, N1373, N1032);
xor XOR2 (N1818, N1812, N197);
not NOT1 (N1819, N1813);
nor NOR4 (N1820, N1819, N462, N1495, N1006);
buf BUF1 (N1821, N1817);
xor XOR2 (N1822, N1816, N288);
buf BUF1 (N1823, N1814);
buf BUF1 (N1824, N1795);
not NOT1 (N1825, N1779);
nor NOR2 (N1826, N1815, N283);
and AND3 (N1827, N1822, N1013, N1577);
or OR3 (N1828, N1825, N657, N403);
buf BUF1 (N1829, N1823);
nand NAND4 (N1830, N1828, N1509, N959, N721);
nor NOR2 (N1831, N1824, N1372);
nand NAND2 (N1832, N1821, N237);
xor XOR2 (N1833, N1827, N294);
xor XOR2 (N1834, N1818, N1747);
nand NAND2 (N1835, N1829, N600);
and AND3 (N1836, N1834, N705, N1559);
or OR2 (N1837, N1807, N299);
nor NOR4 (N1838, N1832, N195, N1315, N1805);
xor XOR2 (N1839, N1836, N1091);
buf BUF1 (N1840, N1803);
buf BUF1 (N1841, N1826);
nor NOR3 (N1842, N1831, N172, N630);
and AND4 (N1843, N1839, N1789, N327, N1730);
and AND3 (N1844, N1838, N620, N690);
nor NOR3 (N1845, N1830, N652, N1646);
and AND3 (N1846, N1844, N1638, N208);
nand NAND4 (N1847, N1843, N1708, N1129, N294);
or OR3 (N1848, N1846, N1207, N385);
buf BUF1 (N1849, N1845);
or OR4 (N1850, N1833, N286, N488, N1028);
buf BUF1 (N1851, N1835);
and AND4 (N1852, N1851, N724, N276, N1810);
and AND2 (N1853, N1842, N1308);
nor NOR4 (N1854, N1850, N1658, N303, N817);
or OR2 (N1855, N1848, N505);
and AND4 (N1856, N1854, N1143, N601, N801);
nand NAND4 (N1857, N1847, N1177, N514, N808);
buf BUF1 (N1858, N1852);
buf BUF1 (N1859, N1856);
and AND4 (N1860, N1858, N1075, N707, N888);
nor NOR2 (N1861, N1855, N1447);
and AND4 (N1862, N1859, N934, N521, N97);
nand NAND2 (N1863, N1853, N670);
and AND3 (N1864, N1841, N604, N1180);
or OR3 (N1865, N1820, N964, N1829);
nor NOR4 (N1866, N1837, N1147, N615, N338);
or OR2 (N1867, N1862, N367);
or OR2 (N1868, N1849, N730);
nand NAND3 (N1869, N1840, N78, N850);
nor NOR2 (N1870, N1863, N1789);
not NOT1 (N1871, N1868);
xor XOR2 (N1872, N1861, N637);
not NOT1 (N1873, N1860);
buf BUF1 (N1874, N1867);
not NOT1 (N1875, N1869);
nor NOR3 (N1876, N1866, N1769, N1001);
and AND2 (N1877, N1864, N546);
or OR3 (N1878, N1874, N1537, N1773);
not NOT1 (N1879, N1876);
and AND3 (N1880, N1857, N658, N1052);
xor XOR2 (N1881, N1879, N1648);
xor XOR2 (N1882, N1870, N923);
buf BUF1 (N1883, N1873);
nor NOR2 (N1884, N1872, N72);
not NOT1 (N1885, N1865);
not NOT1 (N1886, N1878);
nand NAND4 (N1887, N1871, N378, N1102, N442);
xor XOR2 (N1888, N1884, N157);
xor XOR2 (N1889, N1883, N1418);
not NOT1 (N1890, N1880);
nand NAND2 (N1891, N1887, N1119);
not NOT1 (N1892, N1891);
nor NOR4 (N1893, N1890, N470, N847, N523);
not NOT1 (N1894, N1875);
nor NOR4 (N1895, N1886, N568, N888, N1608);
not NOT1 (N1896, N1894);
buf BUF1 (N1897, N1896);
xor XOR2 (N1898, N1897, N624);
xor XOR2 (N1899, N1888, N1272);
xor XOR2 (N1900, N1892, N52);
and AND2 (N1901, N1881, N187);
not NOT1 (N1902, N1885);
xor XOR2 (N1903, N1901, N372);
or OR4 (N1904, N1902, N68, N1192, N1113);
buf BUF1 (N1905, N1899);
buf BUF1 (N1906, N1905);
or OR3 (N1907, N1895, N202, N1089);
not NOT1 (N1908, N1877);
buf BUF1 (N1909, N1904);
not NOT1 (N1910, N1900);
nand NAND3 (N1911, N1906, N71, N54);
not NOT1 (N1912, N1882);
nand NAND4 (N1913, N1910, N1616, N1330, N754);
nand NAND2 (N1914, N1893, N1007);
not NOT1 (N1915, N1909);
nand NAND3 (N1916, N1912, N566, N946);
and AND4 (N1917, N1908, N679, N1655, N1200);
or OR4 (N1918, N1914, N716, N1173, N530);
not NOT1 (N1919, N1913);
buf BUF1 (N1920, N1911);
buf BUF1 (N1921, N1889);
and AND2 (N1922, N1917, N1333);
nand NAND2 (N1923, N1922, N1280);
xor XOR2 (N1924, N1921, N421);
nor NOR4 (N1925, N1923, N1019, N579, N997);
and AND3 (N1926, N1918, N1149, N551);
xor XOR2 (N1927, N1907, N369);
not NOT1 (N1928, N1924);
not NOT1 (N1929, N1903);
nand NAND4 (N1930, N1919, N696, N1191, N545);
not NOT1 (N1931, N1916);
and AND2 (N1932, N1915, N91);
xor XOR2 (N1933, N1928, N403);
buf BUF1 (N1934, N1898);
nand NAND4 (N1935, N1926, N957, N1166, N1842);
and AND3 (N1936, N1925, N468, N1531);
xor XOR2 (N1937, N1930, N1076);
or OR4 (N1938, N1931, N226, N1472, N1440);
nand NAND4 (N1939, N1935, N333, N786, N479);
nand NAND4 (N1940, N1936, N87, N1831, N68);
nor NOR2 (N1941, N1937, N953);
and AND4 (N1942, N1933, N1684, N864, N1810);
buf BUF1 (N1943, N1920);
and AND3 (N1944, N1943, N1730, N1610);
nand NAND2 (N1945, N1940, N1235);
buf BUF1 (N1946, N1932);
not NOT1 (N1947, N1927);
nor NOR4 (N1948, N1929, N1940, N556, N1679);
xor XOR2 (N1949, N1942, N1473);
and AND3 (N1950, N1941, N1563, N982);
and AND3 (N1951, N1947, N904, N608);
nand NAND3 (N1952, N1948, N862, N399);
and AND4 (N1953, N1952, N661, N1481, N926);
buf BUF1 (N1954, N1939);
or OR3 (N1955, N1944, N1080, N525);
and AND3 (N1956, N1949, N1462, N1093);
and AND2 (N1957, N1950, N1483);
and AND2 (N1958, N1956, N453);
nand NAND3 (N1959, N1945, N1170, N394);
and AND2 (N1960, N1957, N786);
nor NOR2 (N1961, N1960, N732);
and AND3 (N1962, N1951, N1560, N846);
nor NOR4 (N1963, N1934, N1836, N1206, N354);
nor NOR3 (N1964, N1963, N7, N543);
buf BUF1 (N1965, N1938);
and AND3 (N1966, N1964, N1152, N1718);
nand NAND2 (N1967, N1955, N1276);
nor NOR4 (N1968, N1959, N1320, N550, N279);
nor NOR3 (N1969, N1946, N961, N1265);
not NOT1 (N1970, N1958);
or OR4 (N1971, N1954, N521, N1232, N740);
or OR4 (N1972, N1970, N1568, N281, N869);
nand NAND4 (N1973, N1971, N1624, N1204, N982);
xor XOR2 (N1974, N1967, N1170);
or OR4 (N1975, N1962, N1032, N461, N141);
and AND2 (N1976, N1966, N1220);
and AND4 (N1977, N1953, N939, N1306, N1062);
xor XOR2 (N1978, N1968, N110);
nor NOR3 (N1979, N1965, N220, N774);
xor XOR2 (N1980, N1979, N658);
not NOT1 (N1981, N1976);
nor NOR2 (N1982, N1961, N1753);
nor NOR3 (N1983, N1974, N99, N538);
and AND3 (N1984, N1982, N850, N1538);
or OR2 (N1985, N1978, N1564);
not NOT1 (N1986, N1985);
and AND3 (N1987, N1975, N233, N1795);
xor XOR2 (N1988, N1984, N1073);
not NOT1 (N1989, N1987);
not NOT1 (N1990, N1989);
xor XOR2 (N1991, N1972, N1506);
xor XOR2 (N1992, N1988, N349);
or OR2 (N1993, N1983, N180);
xor XOR2 (N1994, N1981, N951);
nor NOR3 (N1995, N1994, N583, N1949);
buf BUF1 (N1996, N1991);
nand NAND4 (N1997, N1973, N623, N987, N305);
nor NOR4 (N1998, N1980, N738, N230, N196);
not NOT1 (N1999, N1997);
buf BUF1 (N2000, N1999);
not NOT1 (N2001, N1995);
buf BUF1 (N2002, N1992);
buf BUF1 (N2003, N1996);
not NOT1 (N2004, N1998);
and AND3 (N2005, N1977, N1349, N179);
nand NAND3 (N2006, N1969, N1676, N104);
not NOT1 (N2007, N2001);
buf BUF1 (N2008, N2002);
xor XOR2 (N2009, N2004, N1330);
or OR4 (N2010, N1993, N49, N1097, N1909);
nor NOR2 (N2011, N1990, N1218);
buf BUF1 (N2012, N2009);
buf BUF1 (N2013, N2000);
nor NOR4 (N2014, N2008, N1180, N1291, N431);
or OR3 (N2015, N1986, N1716, N136);
nor NOR4 (N2016, N2010, N1475, N215, N915);
and AND3 (N2017, N2012, N1683, N553);
not NOT1 (N2018, N2017);
and AND3 (N2019, N2006, N587, N1998);
or OR3 (N2020, N2015, N1011, N1105);
not NOT1 (N2021, N2003);
or OR4 (N2022, N2021, N75, N829, N327);
not NOT1 (N2023, N2018);
nand NAND4 (N2024, N2016, N82, N836, N487);
or OR3 (N2025, N2005, N1732, N910);
nand NAND3 (N2026, N2011, N820, N921);
not NOT1 (N2027, N2014);
nor NOR2 (N2028, N2007, N880);
and AND4 (N2029, N2019, N100, N458, N420);
nand NAND2 (N2030, N2013, N1664);
buf BUF1 (N2031, N2020);
and AND3 (N2032, N2029, N1184, N221);
nor NOR4 (N2033, N2028, N672, N915, N1838);
xor XOR2 (N2034, N2027, N1259);
not NOT1 (N2035, N2033);
or OR3 (N2036, N2030, N1074, N127);
not NOT1 (N2037, N2026);
and AND3 (N2038, N2036, N1218, N1107);
and AND3 (N2039, N2031, N1292, N662);
nand NAND2 (N2040, N2039, N68);
or OR2 (N2041, N2038, N1427);
nor NOR2 (N2042, N2024, N528);
buf BUF1 (N2043, N2022);
nand NAND3 (N2044, N2043, N197, N1714);
nand NAND4 (N2045, N2023, N843, N1094, N125);
nor NOR2 (N2046, N2025, N1400);
not NOT1 (N2047, N2044);
xor XOR2 (N2048, N2040, N1118);
buf BUF1 (N2049, N2032);
nand NAND4 (N2050, N2049, N1558, N1834, N302);
or OR3 (N2051, N2035, N1862, N642);
and AND2 (N2052, N2042, N1590);
xor XOR2 (N2053, N2046, N1885);
nand NAND2 (N2054, N2052, N231);
nand NAND4 (N2055, N2050, N719, N242, N1609);
nand NAND2 (N2056, N2037, N192);
not NOT1 (N2057, N2053);
nor NOR3 (N2058, N2056, N1693, N1806);
xor XOR2 (N2059, N2047, N1275);
nand NAND3 (N2060, N2059, N102, N640);
buf BUF1 (N2061, N2041);
not NOT1 (N2062, N2061);
and AND3 (N2063, N2055, N1961, N910);
and AND4 (N2064, N2060, N971, N1607, N784);
and AND2 (N2065, N2058, N1899);
or OR2 (N2066, N2051, N1092);
xor XOR2 (N2067, N2048, N1898);
buf BUF1 (N2068, N2067);
xor XOR2 (N2069, N2062, N567);
buf BUF1 (N2070, N2034);
buf BUF1 (N2071, N2070);
buf BUF1 (N2072, N2054);
buf BUF1 (N2073, N2072);
not NOT1 (N2074, N2065);
nor NOR3 (N2075, N2057, N258, N1927);
nor NOR4 (N2076, N2063, N848, N442, N63);
nor NOR4 (N2077, N2073, N1090, N1275, N1145);
nor NOR4 (N2078, N2076, N1551, N1573, N1765);
and AND4 (N2079, N2068, N1780, N1433, N1770);
nand NAND2 (N2080, N2071, N1594);
nand NAND4 (N2081, N2069, N1646, N443, N983);
buf BUF1 (N2082, N2066);
and AND2 (N2083, N2077, N357);
buf BUF1 (N2084, N2064);
nor NOR4 (N2085, N2080, N606, N810, N1209);
xor XOR2 (N2086, N2045, N736);
nand NAND2 (N2087, N2081, N1537);
nand NAND3 (N2088, N2078, N1324, N1960);
xor XOR2 (N2089, N2074, N1826);
not NOT1 (N2090, N2082);
xor XOR2 (N2091, N2083, N1848);
xor XOR2 (N2092, N2089, N1389);
buf BUF1 (N2093, N2088);
xor XOR2 (N2094, N2090, N2001);
xor XOR2 (N2095, N2079, N1853);
buf BUF1 (N2096, N2087);
nand NAND2 (N2097, N2075, N471);
not NOT1 (N2098, N2092);
buf BUF1 (N2099, N2091);
or OR2 (N2100, N2084, N398);
nand NAND2 (N2101, N2086, N12);
xor XOR2 (N2102, N2085, N1730);
or OR2 (N2103, N2094, N1134);
nand NAND2 (N2104, N2093, N1106);
xor XOR2 (N2105, N2100, N1690);
xor XOR2 (N2106, N2098, N774);
buf BUF1 (N2107, N2095);
xor XOR2 (N2108, N2096, N1648);
and AND2 (N2109, N2106, N1656);
buf BUF1 (N2110, N2105);
nor NOR3 (N2111, N2102, N64, N1874);
nor NOR2 (N2112, N2103, N462);
or OR2 (N2113, N2109, N1900);
or OR4 (N2114, N2110, N1693, N1141, N513);
nand NAND3 (N2115, N2097, N294, N678);
not NOT1 (N2116, N2104);
nand NAND4 (N2117, N2114, N281, N1447, N773);
or OR2 (N2118, N2108, N1734);
nand NAND4 (N2119, N2118, N628, N1051, N43);
and AND4 (N2120, N2107, N1176, N669, N194);
buf BUF1 (N2121, N2112);
nand NAND3 (N2122, N2115, N859, N452);
xor XOR2 (N2123, N2116, N524);
or OR3 (N2124, N2120, N538, N1907);
buf BUF1 (N2125, N2124);
buf BUF1 (N2126, N2123);
nor NOR2 (N2127, N2125, N29);
xor XOR2 (N2128, N2113, N1835);
and AND2 (N2129, N2101, N1360);
not NOT1 (N2130, N2129);
not NOT1 (N2131, N2126);
nor NOR4 (N2132, N2122, N1311, N182, N1436);
and AND3 (N2133, N2130, N2055, N1117);
and AND3 (N2134, N2133, N2064, N1863);
nand NAND2 (N2135, N2134, N1051);
nand NAND4 (N2136, N2119, N1830, N1987, N1557);
or OR2 (N2137, N2136, N2095);
nor NOR4 (N2138, N2111, N1325, N422, N1800);
not NOT1 (N2139, N2138);
and AND3 (N2140, N2137, N454, N1856);
not NOT1 (N2141, N2139);
nor NOR4 (N2142, N2140, N1096, N1176, N1141);
nor NOR2 (N2143, N2128, N2136);
xor XOR2 (N2144, N2142, N1175);
or OR2 (N2145, N2135, N1462);
not NOT1 (N2146, N2099);
and AND3 (N2147, N2131, N922, N2060);
buf BUF1 (N2148, N2132);
xor XOR2 (N2149, N2146, N995);
and AND2 (N2150, N2143, N2137);
nand NAND4 (N2151, N2150, N2114, N904, N42);
nand NAND2 (N2152, N2145, N1782);
nor NOR2 (N2153, N2144, N1348);
or OR3 (N2154, N2153, N1677, N617);
or OR4 (N2155, N2141, N843, N1757, N83);
and AND4 (N2156, N2151, N1966, N1596, N695);
and AND3 (N2157, N2152, N1148, N227);
not NOT1 (N2158, N2117);
buf BUF1 (N2159, N2154);
xor XOR2 (N2160, N2155, N1948);
and AND2 (N2161, N2147, N189);
or OR4 (N2162, N2156, N959, N671, N1435);
not NOT1 (N2163, N2148);
nor NOR4 (N2164, N2121, N1103, N2082, N1287);
or OR2 (N2165, N2161, N460);
and AND3 (N2166, N2158, N755, N472);
not NOT1 (N2167, N2157);
not NOT1 (N2168, N2160);
or OR3 (N2169, N2165, N1413, N700);
buf BUF1 (N2170, N2168);
nand NAND2 (N2171, N2167, N473);
nor NOR2 (N2172, N2162, N855);
xor XOR2 (N2173, N2149, N648);
not NOT1 (N2174, N2170);
xor XOR2 (N2175, N2127, N315);
buf BUF1 (N2176, N2172);
nand NAND4 (N2177, N2166, N1113, N908, N20);
buf BUF1 (N2178, N2171);
or OR4 (N2179, N2164, N494, N2010, N2068);
not NOT1 (N2180, N2177);
nand NAND4 (N2181, N2178, N1349, N1611, N894);
and AND2 (N2182, N2179, N361);
nor NOR4 (N2183, N2159, N982, N602, N103);
nand NAND4 (N2184, N2176, N1477, N1668, N380);
xor XOR2 (N2185, N2182, N577);
not NOT1 (N2186, N2180);
and AND2 (N2187, N2186, N1571);
not NOT1 (N2188, N2181);
buf BUF1 (N2189, N2185);
nand NAND3 (N2190, N2163, N1528, N1891);
or OR4 (N2191, N2184, N593, N1211, N2063);
buf BUF1 (N2192, N2190);
not NOT1 (N2193, N2192);
nand NAND2 (N2194, N2193, N609);
xor XOR2 (N2195, N2187, N674);
not NOT1 (N2196, N2175);
and AND2 (N2197, N2183, N2022);
nor NOR3 (N2198, N2188, N416, N362);
and AND2 (N2199, N2191, N2061);
nor NOR4 (N2200, N2194, N1637, N86, N2106);
or OR3 (N2201, N2173, N1263, N2081);
nand NAND3 (N2202, N2201, N503, N1208);
nand NAND4 (N2203, N2195, N2180, N575, N1181);
and AND2 (N2204, N2202, N1758);
nand NAND4 (N2205, N2200, N528, N1358, N1919);
buf BUF1 (N2206, N2205);
and AND3 (N2207, N2206, N2037, N424);
buf BUF1 (N2208, N2189);
buf BUF1 (N2209, N2203);
or OR3 (N2210, N2198, N1369, N1978);
buf BUF1 (N2211, N2174);
or OR4 (N2212, N2199, N1718, N360, N443);
buf BUF1 (N2213, N2209);
or OR2 (N2214, N2207, N681);
not NOT1 (N2215, N2196);
or OR2 (N2216, N2214, N875);
buf BUF1 (N2217, N2204);
and AND4 (N2218, N2216, N1472, N74, N498);
and AND3 (N2219, N2212, N1710, N1593);
nor NOR3 (N2220, N2218, N1248, N1461);
buf BUF1 (N2221, N2208);
buf BUF1 (N2222, N2210);
not NOT1 (N2223, N2211);
or OR4 (N2224, N2213, N1961, N1138, N1192);
xor XOR2 (N2225, N2223, N1528);
and AND3 (N2226, N2224, N1643, N1296);
not NOT1 (N2227, N2219);
and AND4 (N2228, N2220, N1554, N1648, N211);
or OR3 (N2229, N2197, N1631, N1978);
xor XOR2 (N2230, N2215, N2108);
and AND4 (N2231, N2230, N1531, N171, N1158);
and AND3 (N2232, N2217, N696, N316);
nand NAND3 (N2233, N2169, N1131, N1064);
buf BUF1 (N2234, N2232);
nor NOR2 (N2235, N2231, N1850);
or OR3 (N2236, N2227, N1137, N429);
or OR3 (N2237, N2222, N475, N346);
xor XOR2 (N2238, N2225, N1637);
nor NOR4 (N2239, N2226, N662, N1475, N961);
buf BUF1 (N2240, N2234);
xor XOR2 (N2241, N2240, N924);
or OR4 (N2242, N2241, N1445, N831, N11);
not NOT1 (N2243, N2242);
not NOT1 (N2244, N2228);
nand NAND4 (N2245, N2244, N243, N723, N82);
buf BUF1 (N2246, N2243);
nand NAND4 (N2247, N2235, N809, N1899, N1946);
nand NAND3 (N2248, N2246, N422, N1355);
buf BUF1 (N2249, N2248);
not NOT1 (N2250, N2237);
or OR4 (N2251, N2233, N284, N1275, N67);
xor XOR2 (N2252, N2229, N52);
xor XOR2 (N2253, N2236, N1272);
and AND2 (N2254, N2252, N152);
and AND4 (N2255, N2239, N874, N1438, N315);
and AND3 (N2256, N2249, N437, N2163);
nand NAND3 (N2257, N2250, N2065, N982);
xor XOR2 (N2258, N2256, N1968);
or OR4 (N2259, N2247, N1835, N1945, N1304);
buf BUF1 (N2260, N2253);
buf BUF1 (N2261, N2259);
or OR4 (N2262, N2221, N1520, N145, N810);
not NOT1 (N2263, N2255);
xor XOR2 (N2264, N2263, N1117);
and AND2 (N2265, N2245, N600);
and AND3 (N2266, N2238, N428, N1630);
not NOT1 (N2267, N2260);
nand NAND3 (N2268, N2266, N1914, N1330);
and AND2 (N2269, N2251, N1839);
not NOT1 (N2270, N2262);
not NOT1 (N2271, N2270);
buf BUF1 (N2272, N2271);
and AND4 (N2273, N2254, N1364, N1299, N598);
xor XOR2 (N2274, N2261, N1445);
nor NOR3 (N2275, N2273, N1995, N2023);
and AND4 (N2276, N2264, N1936, N816, N432);
or OR4 (N2277, N2268, N947, N1313, N1280);
buf BUF1 (N2278, N2272);
xor XOR2 (N2279, N2277, N1996);
and AND4 (N2280, N2269, N895, N1501, N1650);
and AND4 (N2281, N2275, N1222, N1204, N953);
xor XOR2 (N2282, N2274, N791);
buf BUF1 (N2283, N2258);
nor NOR4 (N2284, N2280, N94, N1143, N777);
nor NOR3 (N2285, N2278, N1067, N1295);
xor XOR2 (N2286, N2284, N1396);
xor XOR2 (N2287, N2265, N2116);
not NOT1 (N2288, N2285);
xor XOR2 (N2289, N2267, N2226);
not NOT1 (N2290, N2288);
buf BUF1 (N2291, N2279);
and AND3 (N2292, N2283, N340, N98);
nand NAND3 (N2293, N2281, N1185, N551);
not NOT1 (N2294, N2257);
nor NOR2 (N2295, N2276, N715);
not NOT1 (N2296, N2287);
nand NAND3 (N2297, N2293, N287, N751);
buf BUF1 (N2298, N2296);
and AND4 (N2299, N2291, N2147, N795, N1213);
and AND4 (N2300, N2292, N1831, N401, N1794);
nor NOR3 (N2301, N2286, N2265, N1086);
nor NOR4 (N2302, N2300, N324, N1635, N1416);
or OR4 (N2303, N2297, N2042, N2236, N1243);
nor NOR3 (N2304, N2299, N696, N1852);
or OR2 (N2305, N2289, N68);
xor XOR2 (N2306, N2302, N1001);
buf BUF1 (N2307, N2301);
xor XOR2 (N2308, N2304, N1281);
xor XOR2 (N2309, N2294, N1951);
and AND3 (N2310, N2308, N375, N1474);
or OR4 (N2311, N2282, N277, N1117, N1779);
nand NAND2 (N2312, N2309, N480);
buf BUF1 (N2313, N2310);
not NOT1 (N2314, N2307);
buf BUF1 (N2315, N2312);
or OR3 (N2316, N2295, N350, N746);
xor XOR2 (N2317, N2314, N1401);
xor XOR2 (N2318, N2311, N1390);
not NOT1 (N2319, N2318);
xor XOR2 (N2320, N2298, N1848);
buf BUF1 (N2321, N2320);
nor NOR2 (N2322, N2303, N772);
or OR2 (N2323, N2305, N1163);
and AND4 (N2324, N2306, N1369, N1675, N389);
nor NOR2 (N2325, N2319, N636);
or OR4 (N2326, N2316, N287, N542, N1358);
and AND2 (N2327, N2325, N2077);
xor XOR2 (N2328, N2290, N1057);
buf BUF1 (N2329, N2313);
nor NOR4 (N2330, N2329, N332, N747, N386);
nor NOR4 (N2331, N2322, N585, N379, N2275);
not NOT1 (N2332, N2328);
buf BUF1 (N2333, N2315);
buf BUF1 (N2334, N2332);
not NOT1 (N2335, N2331);
nand NAND2 (N2336, N2323, N1034);
xor XOR2 (N2337, N2321, N561);
or OR4 (N2338, N2330, N589, N1827, N1064);
nor NOR2 (N2339, N2333, N68);
not NOT1 (N2340, N2339);
xor XOR2 (N2341, N2335, N1506);
not NOT1 (N2342, N2340);
and AND3 (N2343, N2317, N818, N2174);
nor NOR2 (N2344, N2336, N732);
nand NAND4 (N2345, N2344, N717, N965, N909);
xor XOR2 (N2346, N2338, N1912);
not NOT1 (N2347, N2342);
xor XOR2 (N2348, N2341, N1345);
nand NAND4 (N2349, N2324, N148, N302, N926);
and AND2 (N2350, N2348, N1722);
or OR2 (N2351, N2337, N223);
or OR2 (N2352, N2351, N1532);
xor XOR2 (N2353, N2350, N131);
buf BUF1 (N2354, N2352);
xor XOR2 (N2355, N2354, N1973);
or OR3 (N2356, N2353, N1912, N160);
nor NOR3 (N2357, N2343, N1092, N2068);
and AND3 (N2358, N2345, N962, N156);
or OR2 (N2359, N2346, N789);
nor NOR2 (N2360, N2349, N1335);
not NOT1 (N2361, N2356);
buf BUF1 (N2362, N2327);
and AND4 (N2363, N2347, N484, N1389, N1817);
nand NAND2 (N2364, N2355, N760);
nand NAND4 (N2365, N2361, N364, N359, N2112);
and AND2 (N2366, N2362, N2299);
or OR4 (N2367, N2360, N921, N2246, N359);
buf BUF1 (N2368, N2363);
not NOT1 (N2369, N2368);
nor NOR4 (N2370, N2359, N606, N569, N578);
buf BUF1 (N2371, N2358);
nor NOR4 (N2372, N2366, N1121, N1909, N2187);
not NOT1 (N2373, N2364);
and AND3 (N2374, N2334, N452, N435);
nor NOR4 (N2375, N2369, N1047, N1408, N575);
nand NAND2 (N2376, N2371, N764);
not NOT1 (N2377, N2367);
xor XOR2 (N2378, N2374, N846);
and AND3 (N2379, N2370, N1342, N553);
or OR3 (N2380, N2326, N2046, N18);
and AND2 (N2381, N2377, N644);
xor XOR2 (N2382, N2380, N2228);
buf BUF1 (N2383, N2378);
nand NAND2 (N2384, N2373, N2053);
and AND3 (N2385, N2379, N1528, N1095);
not NOT1 (N2386, N2385);
or OR3 (N2387, N2372, N1831, N697);
nand NAND4 (N2388, N2376, N27, N1800, N463);
buf BUF1 (N2389, N2375);
and AND2 (N2390, N2388, N284);
xor XOR2 (N2391, N2389, N946);
nor NOR4 (N2392, N2365, N991, N1167, N1432);
or OR2 (N2393, N2391, N582);
or OR4 (N2394, N2390, N69, N1079, N1728);
xor XOR2 (N2395, N2392, N1569);
xor XOR2 (N2396, N2381, N2222);
xor XOR2 (N2397, N2394, N1258);
or OR4 (N2398, N2397, N2345, N782, N3);
nor NOR4 (N2399, N2387, N2275, N194, N553);
and AND2 (N2400, N2384, N1163);
xor XOR2 (N2401, N2382, N176);
not NOT1 (N2402, N2401);
nor NOR4 (N2403, N2383, N383, N986, N603);
and AND2 (N2404, N2386, N182);
nor NOR4 (N2405, N2400, N898, N1759, N338);
nor NOR2 (N2406, N2396, N1699);
or OR2 (N2407, N2399, N1222);
nand NAND2 (N2408, N2393, N644);
and AND4 (N2409, N2407, N1368, N146, N24);
xor XOR2 (N2410, N2404, N276);
not NOT1 (N2411, N2409);
nor NOR4 (N2412, N2395, N1541, N1790, N1334);
and AND2 (N2413, N2410, N264);
and AND4 (N2414, N2411, N2072, N837, N1822);
xor XOR2 (N2415, N2412, N1892);
not NOT1 (N2416, N2405);
buf BUF1 (N2417, N2402);
and AND3 (N2418, N2357, N1377, N585);
buf BUF1 (N2419, N2408);
buf BUF1 (N2420, N2406);
not NOT1 (N2421, N2420);
nand NAND4 (N2422, N2418, N1577, N797, N2354);
xor XOR2 (N2423, N2415, N1643);
buf BUF1 (N2424, N2416);
xor XOR2 (N2425, N2422, N2295);
xor XOR2 (N2426, N2413, N414);
or OR3 (N2427, N2425, N1910, N1058);
or OR3 (N2428, N2417, N129, N886);
and AND2 (N2429, N2423, N110);
xor XOR2 (N2430, N2428, N799);
xor XOR2 (N2431, N2430, N219);
buf BUF1 (N2432, N2403);
nand NAND3 (N2433, N2398, N1194, N1754);
buf BUF1 (N2434, N2421);
or OR2 (N2435, N2427, N932);
not NOT1 (N2436, N2434);
xor XOR2 (N2437, N2424, N1177);
xor XOR2 (N2438, N2432, N1816);
or OR4 (N2439, N2436, N357, N992, N26);
and AND2 (N2440, N2429, N574);
nand NAND2 (N2441, N2426, N1731);
nor NOR3 (N2442, N2439, N1515, N1571);
nor NOR3 (N2443, N2414, N1678, N2403);
and AND2 (N2444, N2431, N448);
xor XOR2 (N2445, N2444, N392);
xor XOR2 (N2446, N2433, N2227);
not NOT1 (N2447, N2445);
or OR2 (N2448, N2443, N2166);
buf BUF1 (N2449, N2447);
and AND2 (N2450, N2441, N98);
nand NAND4 (N2451, N2438, N50, N1806, N1800);
buf BUF1 (N2452, N2446);
nor NOR4 (N2453, N2440, N156, N1084, N1132);
or OR4 (N2454, N2419, N2325, N124, N1945);
or OR4 (N2455, N2435, N13, N1835, N373);
nor NOR2 (N2456, N2451, N2206);
or OR4 (N2457, N2437, N432, N2108, N1198);
nand NAND2 (N2458, N2450, N1149);
nor NOR3 (N2459, N2442, N1484, N1288);
nand NAND4 (N2460, N2456, N1535, N367, N2055);
nor NOR2 (N2461, N2458, N1848);
nor NOR4 (N2462, N2454, N624, N541, N771);
not NOT1 (N2463, N2448);
nor NOR3 (N2464, N2457, N1414, N728);
or OR3 (N2465, N2455, N375, N581);
and AND4 (N2466, N2449, N654, N1643, N2044);
buf BUF1 (N2467, N2464);
nor NOR3 (N2468, N2453, N889, N1423);
nor NOR4 (N2469, N2465, N1611, N1115, N72);
xor XOR2 (N2470, N2469, N2006);
nor NOR4 (N2471, N2463, N2289, N690, N2295);
buf BUF1 (N2472, N2461);
or OR3 (N2473, N2468, N2296, N329);
xor XOR2 (N2474, N2452, N1962);
nand NAND3 (N2475, N2472, N122, N2049);
xor XOR2 (N2476, N2470, N1415);
xor XOR2 (N2477, N2467, N79);
nor NOR3 (N2478, N2460, N1171, N102);
or OR3 (N2479, N2459, N2119, N1749);
and AND4 (N2480, N2462, N1158, N672, N1708);
and AND2 (N2481, N2480, N1722);
nor NOR4 (N2482, N2475, N437, N895, N779);
or OR4 (N2483, N2474, N137, N1344, N795);
not NOT1 (N2484, N2482);
not NOT1 (N2485, N2466);
and AND4 (N2486, N2479, N2272, N2420, N395);
xor XOR2 (N2487, N2481, N1083);
not NOT1 (N2488, N2487);
buf BUF1 (N2489, N2483);
or OR3 (N2490, N2478, N380, N613);
nand NAND3 (N2491, N2490, N47, N472);
xor XOR2 (N2492, N2484, N805);
nand NAND4 (N2493, N2471, N52, N46, N1799);
nand NAND4 (N2494, N2491, N1213, N1872, N761);
not NOT1 (N2495, N2485);
nand NAND2 (N2496, N2492, N1943);
buf BUF1 (N2497, N2494);
and AND4 (N2498, N2496, N1851, N1397, N2460);
xor XOR2 (N2499, N2489, N1421);
and AND3 (N2500, N2476, N217, N2490);
and AND3 (N2501, N2500, N2045, N772);
or OR2 (N2502, N2473, N1637);
buf BUF1 (N2503, N2493);
not NOT1 (N2504, N2488);
nor NOR4 (N2505, N2495, N1281, N1043, N1221);
buf BUF1 (N2506, N2504);
nor NOR2 (N2507, N2506, N2430);
nand NAND2 (N2508, N2498, N604);
buf BUF1 (N2509, N2497);
nor NOR2 (N2510, N2502, N1921);
or OR4 (N2511, N2486, N1551, N981, N1254);
xor XOR2 (N2512, N2509, N1071);
xor XOR2 (N2513, N2505, N1651);
and AND3 (N2514, N2477, N1784, N856);
nand NAND2 (N2515, N2514, N546);
xor XOR2 (N2516, N2503, N692);
nand NAND2 (N2517, N2508, N2124);
buf BUF1 (N2518, N2511);
nor NOR4 (N2519, N2515, N1426, N1832, N1398);
and AND2 (N2520, N2501, N643);
or OR3 (N2521, N2516, N408, N1244);
and AND2 (N2522, N2517, N2372);
or OR3 (N2523, N2522, N2474, N1696);
buf BUF1 (N2524, N2520);
xor XOR2 (N2525, N2523, N1755);
and AND2 (N2526, N2524, N1359);
not NOT1 (N2527, N2525);
nor NOR4 (N2528, N2518, N2509, N1416, N2333);
nor NOR4 (N2529, N2527, N1680, N1637, N658);
or OR4 (N2530, N2512, N19, N1885, N2096);
xor XOR2 (N2531, N2510, N608);
and AND2 (N2532, N2531, N64);
and AND3 (N2533, N2513, N1199, N1755);
buf BUF1 (N2534, N2530);
buf BUF1 (N2535, N2499);
buf BUF1 (N2536, N2526);
xor XOR2 (N2537, N2535, N2438);
nand NAND3 (N2538, N2536, N2487, N1307);
buf BUF1 (N2539, N2519);
and AND2 (N2540, N2507, N393);
nand NAND2 (N2541, N2533, N1114);
not NOT1 (N2542, N2534);
buf BUF1 (N2543, N2539);
nor NOR3 (N2544, N2542, N2122, N63);
nand NAND3 (N2545, N2528, N1248, N2075);
and AND3 (N2546, N2545, N850, N441);
xor XOR2 (N2547, N2521, N1180);
not NOT1 (N2548, N2547);
buf BUF1 (N2549, N2543);
nor NOR2 (N2550, N2538, N691);
or OR4 (N2551, N2532, N1619, N1274, N2402);
not NOT1 (N2552, N2551);
or OR2 (N2553, N2552, N271);
nand NAND4 (N2554, N2548, N1515, N978, N1824);
and AND3 (N2555, N2549, N1319, N1371);
buf BUF1 (N2556, N2537);
nand NAND3 (N2557, N2540, N2277, N972);
xor XOR2 (N2558, N2553, N822);
and AND4 (N2559, N2550, N2392, N1007, N166);
nor NOR4 (N2560, N2554, N918, N838, N1327);
nor NOR3 (N2561, N2559, N2132, N1374);
xor XOR2 (N2562, N2557, N2157);
and AND2 (N2563, N2555, N1502);
and AND4 (N2564, N2562, N1627, N123, N1347);
nand NAND4 (N2565, N2556, N322, N1461, N837);
nand NAND4 (N2566, N2563, N2075, N1952, N939);
xor XOR2 (N2567, N2546, N1444);
or OR2 (N2568, N2529, N2504);
nor NOR4 (N2569, N2558, N1074, N1542, N731);
buf BUF1 (N2570, N2560);
buf BUF1 (N2571, N2570);
buf BUF1 (N2572, N2541);
nor NOR4 (N2573, N2564, N645, N514, N2387);
nand NAND2 (N2574, N2565, N2282);
not NOT1 (N2575, N2573);
nor NOR4 (N2576, N2575, N1280, N30, N2247);
xor XOR2 (N2577, N2576, N475);
nand NAND2 (N2578, N2566, N2094);
buf BUF1 (N2579, N2572);
and AND4 (N2580, N2574, N1049, N1421, N57);
or OR4 (N2581, N2579, N989, N1496, N521);
or OR3 (N2582, N2577, N194, N2532);
nor NOR2 (N2583, N2578, N498);
or OR4 (N2584, N2583, N1689, N1828, N2582);
not NOT1 (N2585, N530);
buf BUF1 (N2586, N2569);
and AND4 (N2587, N2581, N1461, N1688, N1308);
or OR4 (N2588, N2571, N1276, N2337, N2161);
not NOT1 (N2589, N2544);
not NOT1 (N2590, N2567);
buf BUF1 (N2591, N2568);
or OR4 (N2592, N2587, N1308, N1526, N1191);
or OR2 (N2593, N2588, N1510);
and AND4 (N2594, N2590, N547, N670, N1424);
nor NOR3 (N2595, N2592, N781, N1427);
or OR2 (N2596, N2589, N1045);
buf BUF1 (N2597, N2586);
nand NAND3 (N2598, N2593, N1572, N1884);
xor XOR2 (N2599, N2597, N2099);
or OR3 (N2600, N2591, N1658, N591);
nor NOR3 (N2601, N2584, N710, N641);
nor NOR3 (N2602, N2595, N2281, N22);
and AND2 (N2603, N2585, N546);
or OR3 (N2604, N2602, N1396, N1484);
buf BUF1 (N2605, N2603);
or OR2 (N2606, N2599, N925);
nor NOR3 (N2607, N2600, N1954, N282);
nand NAND4 (N2608, N2580, N1028, N2408, N1589);
nor NOR3 (N2609, N2607, N1481, N1185);
or OR3 (N2610, N2605, N920, N1737);
nand NAND2 (N2611, N2598, N98);
xor XOR2 (N2612, N2611, N482);
nor NOR3 (N2613, N2609, N79, N160);
nor NOR3 (N2614, N2594, N2487, N2248);
buf BUF1 (N2615, N2606);
and AND2 (N2616, N2614, N734);
or OR4 (N2617, N2608, N717, N1327, N1120);
and AND4 (N2618, N2615, N1930, N1496, N1398);
xor XOR2 (N2619, N2561, N444);
nor NOR2 (N2620, N2612, N2126);
nor NOR4 (N2621, N2610, N2249, N684, N550);
and AND3 (N2622, N2613, N1065, N204);
and AND3 (N2623, N2622, N2442, N1971);
and AND4 (N2624, N2619, N209, N1763, N1965);
xor XOR2 (N2625, N2616, N1740);
xor XOR2 (N2626, N2621, N1388);
nand NAND4 (N2627, N2626, N2252, N131, N746);
buf BUF1 (N2628, N2604);
buf BUF1 (N2629, N2601);
buf BUF1 (N2630, N2628);
not NOT1 (N2631, N2620);
buf BUF1 (N2632, N2630);
not NOT1 (N2633, N2624);
or OR2 (N2634, N2623, N1304);
and AND3 (N2635, N2617, N2377, N104);
and AND2 (N2636, N2631, N2289);
not NOT1 (N2637, N2625);
or OR2 (N2638, N2629, N1423);
buf BUF1 (N2639, N2618);
or OR3 (N2640, N2638, N27, N1882);
buf BUF1 (N2641, N2633);
nor NOR2 (N2642, N2640, N824);
nor NOR2 (N2643, N2636, N830);
not NOT1 (N2644, N2632);
nand NAND3 (N2645, N2635, N2107, N2239);
and AND3 (N2646, N2627, N449, N1071);
xor XOR2 (N2647, N2644, N346);
not NOT1 (N2648, N2647);
nor NOR4 (N2649, N2646, N1402, N2292, N1897);
nor NOR4 (N2650, N2596, N1631, N858, N750);
xor XOR2 (N2651, N2648, N2028);
not NOT1 (N2652, N2634);
nor NOR3 (N2653, N2641, N2253, N1383);
buf BUF1 (N2654, N2642);
not NOT1 (N2655, N2639);
not NOT1 (N2656, N2655);
nor NOR3 (N2657, N2650, N708, N2457);
not NOT1 (N2658, N2656);
xor XOR2 (N2659, N2653, N568);
not NOT1 (N2660, N2659);
or OR2 (N2661, N2651, N1532);
not NOT1 (N2662, N2657);
or OR2 (N2663, N2637, N1966);
buf BUF1 (N2664, N2663);
nand NAND2 (N2665, N2658, N177);
and AND4 (N2666, N2664, N2600, N843, N111);
xor XOR2 (N2667, N2666, N160);
and AND4 (N2668, N2660, N2419, N772, N2544);
or OR2 (N2669, N2643, N1672);
nand NAND2 (N2670, N2668, N285);
xor XOR2 (N2671, N2667, N279);
nor NOR3 (N2672, N2662, N2295, N818);
and AND3 (N2673, N2672, N2054, N2632);
and AND4 (N2674, N2670, N1987, N1985, N1129);
xor XOR2 (N2675, N2645, N1502);
not NOT1 (N2676, N2673);
nand NAND2 (N2677, N2654, N1121);
not NOT1 (N2678, N2649);
and AND3 (N2679, N2661, N1497, N1383);
or OR4 (N2680, N2671, N1973, N937, N2367);
nand NAND4 (N2681, N2677, N1291, N821, N2492);
nor NOR4 (N2682, N2665, N443, N601, N848);
or OR4 (N2683, N2669, N2163, N2457, N1068);
nand NAND4 (N2684, N2681, N869, N574, N2366);
or OR4 (N2685, N2652, N851, N2519, N2329);
nor NOR2 (N2686, N2680, N2508);
and AND4 (N2687, N2676, N2328, N256, N628);
xor XOR2 (N2688, N2678, N1463);
buf BUF1 (N2689, N2685);
or OR4 (N2690, N2684, N41, N2241, N616);
nor NOR3 (N2691, N2690, N766, N1137);
nand NAND3 (N2692, N2674, N2558, N403);
or OR3 (N2693, N2687, N209, N1783);
buf BUF1 (N2694, N2692);
not NOT1 (N2695, N2675);
buf BUF1 (N2696, N2683);
buf BUF1 (N2697, N2688);
not NOT1 (N2698, N2694);
or OR4 (N2699, N2697, N2457, N825, N363);
or OR2 (N2700, N2691, N1464);
nor NOR3 (N2701, N2679, N1705, N2458);
and AND3 (N2702, N2700, N1427, N1857);
nand NAND4 (N2703, N2689, N1163, N263, N2085);
or OR2 (N2704, N2698, N500);
xor XOR2 (N2705, N2693, N104);
buf BUF1 (N2706, N2705);
and AND4 (N2707, N2706, N2281, N1313, N1818);
xor XOR2 (N2708, N2704, N1994);
buf BUF1 (N2709, N2696);
and AND2 (N2710, N2695, N1472);
nand NAND2 (N2711, N2707, N1567);
and AND2 (N2712, N2711, N2167);
or OR3 (N2713, N2703, N1696, N2184);
xor XOR2 (N2714, N2712, N660);
or OR4 (N2715, N2701, N2014, N790, N2450);
or OR2 (N2716, N2699, N1324);
not NOT1 (N2717, N2709);
xor XOR2 (N2718, N2682, N1523);
xor XOR2 (N2719, N2716, N24);
nand NAND3 (N2720, N2686, N2610, N2200);
not NOT1 (N2721, N2713);
nand NAND2 (N2722, N2717, N1799);
buf BUF1 (N2723, N2702);
and AND4 (N2724, N2708, N1504, N220, N1226);
buf BUF1 (N2725, N2719);
nand NAND4 (N2726, N2710, N1858, N272, N1109);
or OR3 (N2727, N2723, N1009, N155);
nor NOR4 (N2728, N2720, N1458, N1481, N1648);
or OR4 (N2729, N2722, N2619, N2316, N122);
nor NOR3 (N2730, N2714, N896, N2494);
and AND3 (N2731, N2727, N1747, N37);
and AND4 (N2732, N2725, N2559, N2516, N2514);
not NOT1 (N2733, N2718);
and AND2 (N2734, N2733, N1448);
nand NAND2 (N2735, N2732, N671);
and AND4 (N2736, N2715, N1443, N425, N1969);
xor XOR2 (N2737, N2729, N18);
nand NAND2 (N2738, N2734, N133);
or OR2 (N2739, N2738, N2411);
and AND4 (N2740, N2726, N1293, N2606, N2231);
not NOT1 (N2741, N2736);
or OR4 (N2742, N2728, N2249, N271, N1853);
or OR3 (N2743, N2735, N448, N324);
and AND3 (N2744, N2741, N1860, N2512);
nor NOR2 (N2745, N2731, N2195);
not NOT1 (N2746, N2730);
not NOT1 (N2747, N2739);
not NOT1 (N2748, N2747);
and AND4 (N2749, N2740, N1681, N1571, N1078);
and AND4 (N2750, N2745, N1686, N1351, N2640);
and AND2 (N2751, N2750, N293);
xor XOR2 (N2752, N2744, N1080);
nand NAND3 (N2753, N2724, N1084, N2523);
and AND3 (N2754, N2752, N256, N793);
nor NOR2 (N2755, N2751, N2077);
xor XOR2 (N2756, N2742, N1382);
and AND2 (N2757, N2753, N2480);
and AND4 (N2758, N2746, N1526, N511, N936);
nand NAND4 (N2759, N2757, N43, N2753, N826);
xor XOR2 (N2760, N2737, N663);
nand NAND2 (N2761, N2756, N129);
nor NOR4 (N2762, N2748, N1508, N2112, N2566);
nand NAND3 (N2763, N2759, N1935, N95);
xor XOR2 (N2764, N2721, N2493);
nor NOR2 (N2765, N2743, N97);
buf BUF1 (N2766, N2758);
or OR3 (N2767, N2754, N1300, N1907);
or OR2 (N2768, N2763, N2485);
buf BUF1 (N2769, N2768);
nand NAND4 (N2770, N2761, N1474, N894, N2116);
and AND2 (N2771, N2749, N2319);
buf BUF1 (N2772, N2767);
nand NAND3 (N2773, N2769, N1707, N2594);
not NOT1 (N2774, N2765);
xor XOR2 (N2775, N2772, N1219);
xor XOR2 (N2776, N2774, N2600);
nor NOR2 (N2777, N2755, N425);
nor NOR3 (N2778, N2776, N1129, N447);
nor NOR3 (N2779, N2762, N311, N1513);
or OR4 (N2780, N2766, N357, N2001, N1912);
nand NAND2 (N2781, N2770, N2607);
nand NAND4 (N2782, N2760, N2210, N135, N155);
or OR3 (N2783, N2781, N1827, N1580);
and AND2 (N2784, N2771, N968);
buf BUF1 (N2785, N2775);
nand NAND3 (N2786, N2782, N1587, N1870);
nor NOR2 (N2787, N2777, N797);
buf BUF1 (N2788, N2785);
and AND4 (N2789, N2786, N912, N1219, N1043);
or OR3 (N2790, N2779, N1093, N2507);
xor XOR2 (N2791, N2788, N307);
xor XOR2 (N2792, N2764, N777);
or OR4 (N2793, N2784, N593, N481, N1991);
and AND4 (N2794, N2773, N1919, N2481, N849);
buf BUF1 (N2795, N2787);
and AND2 (N2796, N2789, N1703);
or OR2 (N2797, N2790, N658);
and AND3 (N2798, N2780, N544, N2383);
xor XOR2 (N2799, N2791, N214);
nor NOR2 (N2800, N2794, N2349);
and AND2 (N2801, N2796, N2118);
or OR3 (N2802, N2792, N1175, N2116);
xor XOR2 (N2803, N2802, N1502);
buf BUF1 (N2804, N2793);
or OR2 (N2805, N2801, N1790);
buf BUF1 (N2806, N2799);
nand NAND4 (N2807, N2804, N405, N1830, N382);
nand NAND4 (N2808, N2803, N2200, N1340, N2450);
nor NOR2 (N2809, N2805, N171);
xor XOR2 (N2810, N2798, N1975);
nor NOR4 (N2811, N2807, N1469, N699, N1537);
buf BUF1 (N2812, N2795);
buf BUF1 (N2813, N2811);
and AND4 (N2814, N2797, N1569, N356, N448);
or OR4 (N2815, N2778, N1685, N1979, N1194);
or OR2 (N2816, N2813, N2110);
buf BUF1 (N2817, N2810);
not NOT1 (N2818, N2806);
not NOT1 (N2819, N2816);
buf BUF1 (N2820, N2817);
nand NAND4 (N2821, N2814, N856, N2183, N2182);
or OR2 (N2822, N2808, N196);
nand NAND4 (N2823, N2822, N105, N453, N2003);
buf BUF1 (N2824, N2800);
not NOT1 (N2825, N2809);
and AND4 (N2826, N2819, N2523, N2442, N1566);
or OR2 (N2827, N2825, N438);
xor XOR2 (N2828, N2824, N2795);
nand NAND2 (N2829, N2828, N1733);
nor NOR4 (N2830, N2827, N2288, N1324, N2455);
nor NOR3 (N2831, N2812, N2117, N558);
xor XOR2 (N2832, N2826, N2210);
buf BUF1 (N2833, N2783);
buf BUF1 (N2834, N2820);
not NOT1 (N2835, N2830);
nand NAND4 (N2836, N2834, N1978, N2190, N2579);
xor XOR2 (N2837, N2836, N2596);
buf BUF1 (N2838, N2837);
buf BUF1 (N2839, N2835);
and AND3 (N2840, N2821, N340, N830);
not NOT1 (N2841, N2818);
buf BUF1 (N2842, N2840);
and AND4 (N2843, N2833, N2762, N61, N2835);
not NOT1 (N2844, N2839);
nor NOR4 (N2845, N2829, N1592, N2026, N2771);
xor XOR2 (N2846, N2844, N426);
xor XOR2 (N2847, N2843, N2393);
buf BUF1 (N2848, N2838);
xor XOR2 (N2849, N2848, N1916);
buf BUF1 (N2850, N2823);
and AND2 (N2851, N2845, N2302);
xor XOR2 (N2852, N2842, N2564);
nor NOR2 (N2853, N2847, N1291);
xor XOR2 (N2854, N2850, N2688);
xor XOR2 (N2855, N2846, N607);
nand NAND2 (N2856, N2849, N173);
or OR2 (N2857, N2853, N2623);
not NOT1 (N2858, N2815);
xor XOR2 (N2859, N2831, N683);
not NOT1 (N2860, N2858);
or OR4 (N2861, N2855, N2313, N7, N1926);
nor NOR2 (N2862, N2857, N1406);
nor NOR4 (N2863, N2852, N747, N238, N291);
xor XOR2 (N2864, N2854, N7);
not NOT1 (N2865, N2856);
or OR4 (N2866, N2860, N2364, N1635, N1277);
buf BUF1 (N2867, N2865);
nand NAND2 (N2868, N2851, N2320);
and AND3 (N2869, N2863, N700, N860);
or OR3 (N2870, N2867, N2045, N168);
not NOT1 (N2871, N2866);
not NOT1 (N2872, N2859);
nand NAND2 (N2873, N2871, N1976);
buf BUF1 (N2874, N2861);
nand NAND3 (N2875, N2869, N2516, N2548);
xor XOR2 (N2876, N2832, N1223);
not NOT1 (N2877, N2870);
nor NOR4 (N2878, N2841, N594, N1198, N578);
and AND2 (N2879, N2876, N1660);
nand NAND4 (N2880, N2877, N402, N2709, N771);
or OR4 (N2881, N2875, N1295, N285, N2231);
or OR2 (N2882, N2879, N900);
or OR3 (N2883, N2873, N285, N798);
nand NAND2 (N2884, N2868, N1565);
not NOT1 (N2885, N2874);
xor XOR2 (N2886, N2864, N2035);
nand NAND4 (N2887, N2881, N2603, N2206, N1895);
buf BUF1 (N2888, N2883);
nor NOR4 (N2889, N2888, N1471, N433, N519);
and AND3 (N2890, N2889, N1400, N1509);
and AND2 (N2891, N2882, N1753);
not NOT1 (N2892, N2872);
and AND3 (N2893, N2890, N63, N2674);
and AND2 (N2894, N2884, N2802);
or OR4 (N2895, N2892, N2868, N110, N1881);
nor NOR3 (N2896, N2895, N1299, N1105);
nor NOR3 (N2897, N2893, N44, N1690);
nor NOR3 (N2898, N2862, N276, N1574);
or OR2 (N2899, N2885, N2320);
buf BUF1 (N2900, N2897);
not NOT1 (N2901, N2898);
xor XOR2 (N2902, N2900, N432);
buf BUF1 (N2903, N2880);
nor NOR4 (N2904, N2899, N135, N741, N850);
and AND2 (N2905, N2902, N1493);
or OR2 (N2906, N2891, N2155);
xor XOR2 (N2907, N2878, N354);
not NOT1 (N2908, N2904);
nor NOR3 (N2909, N2903, N992, N2367);
or OR2 (N2910, N2894, N93);
or OR2 (N2911, N2905, N1572);
and AND3 (N2912, N2896, N887, N1520);
xor XOR2 (N2913, N2911, N42);
not NOT1 (N2914, N2908);
and AND3 (N2915, N2906, N1082, N537);
or OR2 (N2916, N2915, N261);
nand NAND2 (N2917, N2907, N2382);
xor XOR2 (N2918, N2887, N2789);
or OR3 (N2919, N2909, N639, N1965);
nor NOR2 (N2920, N2917, N990);
and AND4 (N2921, N2886, N1568, N1698, N1522);
and AND2 (N2922, N2912, N323);
not NOT1 (N2923, N2920);
nor NOR2 (N2924, N2923, N908);
xor XOR2 (N2925, N2914, N2827);
or OR2 (N2926, N2901, N1846);
and AND4 (N2927, N2921, N2498, N1677, N349);
and AND2 (N2928, N2927, N1765);
nor NOR2 (N2929, N2919, N180);
not NOT1 (N2930, N2926);
not NOT1 (N2931, N2930);
xor XOR2 (N2932, N2925, N2585);
nand NAND2 (N2933, N2922, N934);
xor XOR2 (N2934, N2928, N2025);
nand NAND4 (N2935, N2933, N667, N864, N2918);
nand NAND3 (N2936, N1214, N1455, N2153);
and AND4 (N2937, N2924, N1916, N2537, N779);
buf BUF1 (N2938, N2931);
and AND4 (N2939, N2929, N1641, N256, N1608);
nor NOR3 (N2940, N2916, N2870, N99);
nand NAND3 (N2941, N2910, N2055, N2181);
xor XOR2 (N2942, N2932, N1364);
buf BUF1 (N2943, N2934);
xor XOR2 (N2944, N2941, N699);
or OR2 (N2945, N2944, N657);
buf BUF1 (N2946, N2939);
and AND4 (N2947, N2940, N2030, N245, N1576);
nor NOR4 (N2948, N2942, N2141, N856, N754);
nor NOR4 (N2949, N2936, N2533, N2020, N2158);
and AND4 (N2950, N2937, N1239, N1180, N1560);
xor XOR2 (N2951, N2948, N944);
or OR3 (N2952, N2943, N1832, N2911);
buf BUF1 (N2953, N2951);
xor XOR2 (N2954, N2947, N1482);
not NOT1 (N2955, N2949);
xor XOR2 (N2956, N2952, N2873);
nand NAND4 (N2957, N2946, N1729, N2250, N2539);
not NOT1 (N2958, N2954);
and AND2 (N2959, N2913, N1022);
and AND4 (N2960, N2950, N56, N63, N54);
not NOT1 (N2961, N2938);
nor NOR4 (N2962, N2957, N2888, N1081, N1201);
and AND2 (N2963, N2958, N1071);
and AND4 (N2964, N2945, N157, N528, N1202);
buf BUF1 (N2965, N2960);
nand NAND3 (N2966, N2963, N2312, N2608);
nor NOR3 (N2967, N2935, N404, N2807);
not NOT1 (N2968, N2962);
and AND4 (N2969, N2968, N466, N2534, N2094);
xor XOR2 (N2970, N2953, N691);
xor XOR2 (N2971, N2959, N572);
nand NAND4 (N2972, N2969, N2519, N395, N283);
and AND2 (N2973, N2965, N1338);
nor NOR4 (N2974, N2961, N2168, N2921, N1302);
nor NOR3 (N2975, N2973, N2354, N2075);
and AND2 (N2976, N2967, N2053);
not NOT1 (N2977, N2972);
nor NOR2 (N2978, N2964, N931);
and AND3 (N2979, N2978, N1963, N2020);
nand NAND4 (N2980, N2974, N1233, N776, N2368);
nand NAND2 (N2981, N2956, N1411);
nor NOR2 (N2982, N2980, N2236);
nand NAND4 (N2983, N2975, N2514, N608, N2354);
buf BUF1 (N2984, N2983);
xor XOR2 (N2985, N2984, N996);
not NOT1 (N2986, N2976);
nor NOR4 (N2987, N2979, N2017, N691, N2019);
buf BUF1 (N2988, N2955);
buf BUF1 (N2989, N2971);
nand NAND3 (N2990, N2966, N1601, N2036);
and AND2 (N2991, N2989, N293);
and AND3 (N2992, N2982, N146, N2492);
xor XOR2 (N2993, N2981, N2060);
or OR3 (N2994, N2987, N1519, N1327);
not NOT1 (N2995, N2990);
nand NAND3 (N2996, N2995, N1351, N2107);
buf BUF1 (N2997, N2996);
nand NAND3 (N2998, N2985, N14, N2473);
nand NAND4 (N2999, N2977, N2856, N2303, N2478);
and AND3 (N3000, N2994, N379, N1791);
or OR2 (N3001, N2986, N516);
and AND3 (N3002, N2970, N1031, N1562);
nor NOR3 (N3003, N2998, N2744, N1476);
and AND4 (N3004, N2993, N1026, N1985, N982);
nand NAND2 (N3005, N2988, N2631);
nor NOR4 (N3006, N3002, N2794, N251, N2149);
or OR3 (N3007, N3005, N1705, N730);
nand NAND4 (N3008, N3003, N1656, N859, N483);
nor NOR3 (N3009, N3006, N2698, N2975);
buf BUF1 (N3010, N3004);
buf BUF1 (N3011, N2999);
or OR2 (N3012, N3000, N2147);
nand NAND2 (N3013, N3010, N2824);
and AND3 (N3014, N3008, N2229, N2835);
not NOT1 (N3015, N3013);
nor NOR2 (N3016, N2997, N1223);
or OR4 (N3017, N3012, N1173, N1977, N1682);
and AND3 (N3018, N3007, N350, N2436);
nand NAND4 (N3019, N3001, N2248, N371, N365);
not NOT1 (N3020, N2991);
xor XOR2 (N3021, N3014, N237);
and AND2 (N3022, N3015, N2195);
not NOT1 (N3023, N3018);
or OR2 (N3024, N3021, N2596);
xor XOR2 (N3025, N2992, N2539);
buf BUF1 (N3026, N3022);
or OR3 (N3027, N3017, N1851, N2886);
nor NOR4 (N3028, N3024, N1109, N1406, N8);
nor NOR4 (N3029, N3009, N2256, N2661, N933);
nand NAND3 (N3030, N3011, N2883, N242);
xor XOR2 (N3031, N3028, N569);
or OR4 (N3032, N3016, N455, N686, N1065);
buf BUF1 (N3033, N3032);
nand NAND2 (N3034, N3029, N981);
and AND3 (N3035, N3023, N1099, N15);
nand NAND4 (N3036, N3020, N1615, N2846, N1395);
nand NAND2 (N3037, N3031, N3014);
nor NOR2 (N3038, N3030, N1766);
nand NAND4 (N3039, N3038, N2110, N938, N2077);
and AND4 (N3040, N3034, N2523, N1668, N2325);
nand NAND4 (N3041, N3035, N2183, N786, N1830);
or OR3 (N3042, N3019, N757, N1485);
buf BUF1 (N3043, N3042);
xor XOR2 (N3044, N3033, N1988);
nor NOR3 (N3045, N3044, N622, N2638);
nand NAND2 (N3046, N3036, N459);
xor XOR2 (N3047, N3026, N5);
buf BUF1 (N3048, N3045);
nand NAND4 (N3049, N3037, N1941, N2486, N492);
nor NOR3 (N3050, N3041, N3036, N2701);
nor NOR3 (N3051, N3043, N915, N1914);
or OR4 (N3052, N3027, N651, N1452, N2467);
not NOT1 (N3053, N3049);
and AND4 (N3054, N3039, N1303, N1242, N1566);
and AND4 (N3055, N3040, N1900, N1603, N2746);
nand NAND3 (N3056, N3051, N2697, N160);
buf BUF1 (N3057, N3056);
and AND3 (N3058, N3053, N2234, N59);
nor NOR2 (N3059, N3054, N1416);
nand NAND3 (N3060, N3058, N2352, N2321);
xor XOR2 (N3061, N3057, N220);
nor NOR3 (N3062, N3047, N2129, N569);
nor NOR3 (N3063, N3062, N118, N2491);
nand NAND4 (N3064, N3055, N2963, N813, N1696);
xor XOR2 (N3065, N3046, N2442);
buf BUF1 (N3066, N3059);
or OR3 (N3067, N3061, N1916, N1375);
nor NOR2 (N3068, N3048, N689);
nor NOR2 (N3069, N3060, N1388);
buf BUF1 (N3070, N3065);
xor XOR2 (N3071, N3069, N1256);
nand NAND4 (N3072, N3025, N826, N2267, N423);
buf BUF1 (N3073, N3063);
buf BUF1 (N3074, N3067);
buf BUF1 (N3075, N3073);
buf BUF1 (N3076, N3074);
buf BUF1 (N3077, N3071);
nand NAND3 (N3078, N3070, N2102, N2628);
not NOT1 (N3079, N3072);
not NOT1 (N3080, N3050);
nand NAND2 (N3081, N3080, N2072);
not NOT1 (N3082, N3068);
or OR2 (N3083, N3079, N1981);
nand NAND4 (N3084, N3075, N1737, N390, N2853);
xor XOR2 (N3085, N3077, N1727);
not NOT1 (N3086, N3083);
xor XOR2 (N3087, N3086, N1734);
and AND4 (N3088, N3081, N1711, N2595, N2178);
nand NAND2 (N3089, N3078, N2867);
not NOT1 (N3090, N3089);
xor XOR2 (N3091, N3084, N2642);
not NOT1 (N3092, N3064);
xor XOR2 (N3093, N3090, N2702);
and AND2 (N3094, N3091, N168);
and AND4 (N3095, N3087, N791, N2427, N553);
xor XOR2 (N3096, N3052, N1035);
not NOT1 (N3097, N3076);
xor XOR2 (N3098, N3085, N1476);
nor NOR3 (N3099, N3092, N682, N2080);
xor XOR2 (N3100, N3093, N166);
or OR4 (N3101, N3097, N536, N268, N1057);
or OR3 (N3102, N3066, N2104, N2796);
buf BUF1 (N3103, N3088);
or OR4 (N3104, N3098, N2264, N266, N1892);
nand NAND2 (N3105, N3103, N609);
nor NOR4 (N3106, N3096, N388, N1458, N2533);
xor XOR2 (N3107, N3095, N464);
xor XOR2 (N3108, N3100, N107);
or OR4 (N3109, N3107, N2201, N661, N2121);
nor NOR4 (N3110, N3102, N1762, N2788, N804);
and AND2 (N3111, N3109, N96);
nand NAND2 (N3112, N3110, N2916);
xor XOR2 (N3113, N3099, N1688);
nand NAND4 (N3114, N3113, N2676, N210, N2781);
xor XOR2 (N3115, N3106, N378);
or OR2 (N3116, N3115, N72);
nor NOR2 (N3117, N3116, N1072);
nand NAND2 (N3118, N3111, N2372);
buf BUF1 (N3119, N3094);
and AND4 (N3120, N3101, N1214, N1199, N2924);
xor XOR2 (N3121, N3114, N1524);
nor NOR3 (N3122, N3082, N2919, N1477);
and AND3 (N3123, N3104, N2939, N2653);
xor XOR2 (N3124, N3112, N2541);
buf BUF1 (N3125, N3121);
or OR2 (N3126, N3122, N1912);
or OR2 (N3127, N3120, N2497);
and AND2 (N3128, N3125, N90);
and AND4 (N3129, N3126, N3009, N2650, N18);
not NOT1 (N3130, N3129);
xor XOR2 (N3131, N3117, N1873);
nand NAND4 (N3132, N3124, N611, N2030, N2276);
or OR4 (N3133, N3127, N1720, N533, N2246);
and AND2 (N3134, N3128, N1977);
or OR2 (N3135, N3108, N2819);
not NOT1 (N3136, N3105);
nand NAND2 (N3137, N3132, N386);
not NOT1 (N3138, N3136);
not NOT1 (N3139, N3123);
or OR3 (N3140, N3119, N941, N1645);
buf BUF1 (N3141, N3139);
buf BUF1 (N3142, N3133);
xor XOR2 (N3143, N3118, N2740);
nor NOR3 (N3144, N3143, N881, N125);
buf BUF1 (N3145, N3137);
and AND3 (N3146, N3134, N1160, N949);
xor XOR2 (N3147, N3141, N1244);
nand NAND3 (N3148, N3145, N318, N339);
xor XOR2 (N3149, N3140, N2113);
nor NOR4 (N3150, N3130, N1538, N1693, N1352);
nor NOR3 (N3151, N3131, N1945, N2437);
or OR4 (N3152, N3146, N2204, N2483, N2330);
buf BUF1 (N3153, N3148);
or OR3 (N3154, N3142, N490, N1226);
nand NAND3 (N3155, N3147, N2587, N1162);
and AND3 (N3156, N3144, N1327, N2140);
buf BUF1 (N3157, N3154);
or OR2 (N3158, N3152, N267);
or OR4 (N3159, N3155, N712, N430, N1343);
and AND3 (N3160, N3153, N100, N2990);
xor XOR2 (N3161, N3157, N885);
nand NAND2 (N3162, N3161, N528);
xor XOR2 (N3163, N3138, N1109);
nor NOR3 (N3164, N3159, N317, N2816);
and AND2 (N3165, N3151, N560);
not NOT1 (N3166, N3149);
nand NAND3 (N3167, N3162, N1134, N773);
xor XOR2 (N3168, N3165, N2427);
nor NOR3 (N3169, N3135, N371, N301);
buf BUF1 (N3170, N3158);
nor NOR4 (N3171, N3169, N1036, N2241, N722);
nor NOR3 (N3172, N3171, N280, N2144);
buf BUF1 (N3173, N3167);
xor XOR2 (N3174, N3173, N2240);
or OR4 (N3175, N3172, N2544, N812, N1419);
buf BUF1 (N3176, N3150);
xor XOR2 (N3177, N3170, N388);
buf BUF1 (N3178, N3160);
buf BUF1 (N3179, N3166);
nor NOR3 (N3180, N3164, N3023, N2222);
not NOT1 (N3181, N3179);
nor NOR4 (N3182, N3168, N1187, N1731, N1201);
and AND4 (N3183, N3175, N784, N742, N1537);
not NOT1 (N3184, N3176);
nor NOR3 (N3185, N3174, N929, N181);
buf BUF1 (N3186, N3178);
not NOT1 (N3187, N3163);
not NOT1 (N3188, N3156);
or OR2 (N3189, N3183, N2047);
not NOT1 (N3190, N3180);
nand NAND4 (N3191, N3181, N334, N1475, N2129);
nand NAND3 (N3192, N3182, N1804, N2092);
buf BUF1 (N3193, N3188);
not NOT1 (N3194, N3184);
or OR2 (N3195, N3189, N2803);
nor NOR4 (N3196, N3185, N2533, N2885, N1454);
xor XOR2 (N3197, N3187, N2413);
and AND3 (N3198, N3196, N892, N328);
nor NOR4 (N3199, N3194, N1876, N2972, N1764);
and AND2 (N3200, N3197, N942);
nand NAND2 (N3201, N3199, N651);
buf BUF1 (N3202, N3198);
buf BUF1 (N3203, N3195);
xor XOR2 (N3204, N3193, N1124);
not NOT1 (N3205, N3191);
or OR2 (N3206, N3192, N2300);
nor NOR4 (N3207, N3204, N572, N923, N865);
buf BUF1 (N3208, N3207);
nor NOR4 (N3209, N3208, N3182, N1997, N1439);
nor NOR4 (N3210, N3201, N876, N508, N47);
nor NOR4 (N3211, N3202, N3144, N1580, N770);
nand NAND3 (N3212, N3210, N1376, N2585);
and AND2 (N3213, N3206, N867);
xor XOR2 (N3214, N3211, N1078);
nor NOR2 (N3215, N3205, N186);
and AND3 (N3216, N3203, N1211, N2342);
not NOT1 (N3217, N3200);
and AND4 (N3218, N3186, N355, N1537, N3196);
buf BUF1 (N3219, N3177);
buf BUF1 (N3220, N3214);
not NOT1 (N3221, N3219);
not NOT1 (N3222, N3209);
or OR3 (N3223, N3190, N900, N647);
buf BUF1 (N3224, N3222);
nand NAND2 (N3225, N3212, N1337);
and AND4 (N3226, N3224, N1512, N863, N1795);
nand NAND2 (N3227, N3225, N1153);
nand NAND3 (N3228, N3221, N871, N2344);
xor XOR2 (N3229, N3217, N2295);
and AND4 (N3230, N3228, N1331, N1589, N1080);
buf BUF1 (N3231, N3230);
buf BUF1 (N3232, N3218);
buf BUF1 (N3233, N3220);
nand NAND3 (N3234, N3226, N1023, N1924);
or OR4 (N3235, N3216, N1605, N2035, N3114);
nand NAND4 (N3236, N3213, N1857, N468, N726);
or OR2 (N3237, N3231, N239);
nor NOR4 (N3238, N3236, N2632, N2679, N586);
or OR4 (N3239, N3238, N2143, N1735, N48);
not NOT1 (N3240, N3234);
or OR3 (N3241, N3227, N597, N682);
nor NOR3 (N3242, N3229, N549, N394);
or OR2 (N3243, N3237, N1821);
or OR4 (N3244, N3241, N1026, N2969, N3107);
xor XOR2 (N3245, N3243, N1957);
and AND3 (N3246, N3223, N2556, N2831);
xor XOR2 (N3247, N3235, N2023);
buf BUF1 (N3248, N3246);
and AND2 (N3249, N3248, N2586);
buf BUF1 (N3250, N3215);
not NOT1 (N3251, N3249);
nor NOR2 (N3252, N3251, N3004);
not NOT1 (N3253, N3247);
and AND4 (N3254, N3245, N1308, N1143, N2747);
nand NAND4 (N3255, N3233, N702, N2393, N2791);
xor XOR2 (N3256, N3242, N606);
and AND2 (N3257, N3253, N2082);
buf BUF1 (N3258, N3244);
or OR3 (N3259, N3240, N855, N1937);
not NOT1 (N3260, N3257);
nand NAND2 (N3261, N3260, N2045);
not NOT1 (N3262, N3258);
nand NAND2 (N3263, N3261, N1071);
not NOT1 (N3264, N3262);
or OR4 (N3265, N3256, N1364, N2367, N2569);
and AND3 (N3266, N3264, N1082, N229);
buf BUF1 (N3267, N3265);
xor XOR2 (N3268, N3259, N1076);
and AND3 (N3269, N3232, N1365, N231);
not NOT1 (N3270, N3269);
buf BUF1 (N3271, N3250);
not NOT1 (N3272, N3252);
and AND3 (N3273, N3271, N1343, N350);
nand NAND4 (N3274, N3267, N1063, N2883, N985);
or OR3 (N3275, N3274, N2129, N924);
xor XOR2 (N3276, N3273, N1982);
and AND2 (N3277, N3239, N180);
and AND3 (N3278, N3266, N2421, N543);
nor NOR3 (N3279, N3278, N2561, N1077);
buf BUF1 (N3280, N3272);
nor NOR2 (N3281, N3268, N281);
nand NAND2 (N3282, N3276, N2086);
not NOT1 (N3283, N3282);
xor XOR2 (N3284, N3280, N2005);
not NOT1 (N3285, N3279);
not NOT1 (N3286, N3283);
xor XOR2 (N3287, N3277, N2665);
nand NAND2 (N3288, N3275, N2418);
nand NAND3 (N3289, N3270, N2787, N2265);
buf BUF1 (N3290, N3281);
nor NOR2 (N3291, N3287, N1096);
buf BUF1 (N3292, N3284);
xor XOR2 (N3293, N3289, N78);
nor NOR4 (N3294, N3263, N881, N2354, N1349);
buf BUF1 (N3295, N3254);
nand NAND3 (N3296, N3290, N225, N2081);
and AND4 (N3297, N3293, N1333, N1932, N2516);
and AND4 (N3298, N3286, N2891, N803, N1182);
nand NAND3 (N3299, N3297, N2756, N2849);
xor XOR2 (N3300, N3296, N2317);
or OR3 (N3301, N3291, N145, N2197);
xor XOR2 (N3302, N3295, N591);
nor NOR3 (N3303, N3302, N1123, N1563);
or OR3 (N3304, N3292, N1424, N1525);
buf BUF1 (N3305, N3301);
not NOT1 (N3306, N3299);
or OR4 (N3307, N3306, N982, N1051, N2661);
and AND3 (N3308, N3288, N1151, N555);
nand NAND4 (N3309, N3298, N2122, N473, N3127);
not NOT1 (N3310, N3255);
nor NOR3 (N3311, N3300, N178, N1783);
nand NAND2 (N3312, N3294, N2295);
not NOT1 (N3313, N3304);
nor NOR2 (N3314, N3305, N658);
nor NOR4 (N3315, N3313, N500, N338, N3118);
or OR3 (N3316, N3315, N2761, N920);
and AND4 (N3317, N3316, N2590, N2750, N150);
and AND4 (N3318, N3303, N2226, N1811, N2917);
nand NAND2 (N3319, N3312, N2719);
not NOT1 (N3320, N3314);
not NOT1 (N3321, N3320);
and AND4 (N3322, N3307, N2728, N2073, N485);
nand NAND2 (N3323, N3317, N1776);
buf BUF1 (N3324, N3321);
xor XOR2 (N3325, N3322, N3166);
buf BUF1 (N3326, N3310);
buf BUF1 (N3327, N3309);
xor XOR2 (N3328, N3319, N1042);
xor XOR2 (N3329, N3311, N1104);
buf BUF1 (N3330, N3328);
nand NAND3 (N3331, N3324, N1239, N175);
or OR4 (N3332, N3330, N1048, N2824, N1141);
nand NAND2 (N3333, N3285, N1765);
nor NOR4 (N3334, N3331, N2147, N253, N1477);
nand NAND3 (N3335, N3327, N2499, N1568);
not NOT1 (N3336, N3333);
xor XOR2 (N3337, N3329, N2602);
buf BUF1 (N3338, N3337);
and AND4 (N3339, N3323, N2028, N1215, N142);
nand NAND3 (N3340, N3308, N3128, N2696);
nor NOR3 (N3341, N3326, N1078, N1867);
buf BUF1 (N3342, N3336);
or OR4 (N3343, N3334, N647, N2354, N152);
buf BUF1 (N3344, N3341);
and AND4 (N3345, N3318, N1824, N3139, N2818);
not NOT1 (N3346, N3332);
nor NOR2 (N3347, N3339, N3031);
xor XOR2 (N3348, N3338, N3086);
nand NAND4 (N3349, N3335, N2627, N653, N1317);
not NOT1 (N3350, N3348);
buf BUF1 (N3351, N3343);
xor XOR2 (N3352, N3325, N2733);
not NOT1 (N3353, N3342);
not NOT1 (N3354, N3351);
or OR3 (N3355, N3345, N2345, N3149);
or OR4 (N3356, N3355, N3129, N658, N1037);
or OR4 (N3357, N3354, N560, N1616, N1542);
nor NOR3 (N3358, N3356, N303, N1310);
nand NAND3 (N3359, N3350, N346, N2641);
buf BUF1 (N3360, N3346);
and AND2 (N3361, N3352, N2788);
nand NAND2 (N3362, N3349, N2901);
or OR3 (N3363, N3362, N2788, N2527);
buf BUF1 (N3364, N3347);
buf BUF1 (N3365, N3340);
nor NOR4 (N3366, N3360, N859, N1043, N2365);
nor NOR2 (N3367, N3361, N3276);
nand NAND4 (N3368, N3353, N583, N2245, N824);
buf BUF1 (N3369, N3365);
or OR3 (N3370, N3367, N2444, N2558);
and AND2 (N3371, N3368, N1846);
or OR2 (N3372, N3369, N3062);
buf BUF1 (N3373, N3366);
buf BUF1 (N3374, N3373);
not NOT1 (N3375, N3364);
or OR3 (N3376, N3363, N261, N2385);
or OR2 (N3377, N3344, N995);
not NOT1 (N3378, N3370);
and AND2 (N3379, N3357, N19);
xor XOR2 (N3380, N3379, N3315);
nor NOR2 (N3381, N3375, N775);
or OR2 (N3382, N3374, N421);
buf BUF1 (N3383, N3377);
nand NAND4 (N3384, N3378, N3104, N723, N3226);
xor XOR2 (N3385, N3358, N2667);
nor NOR4 (N3386, N3380, N1134, N3100, N244);
nor NOR3 (N3387, N3371, N734, N2480);
nor NOR4 (N3388, N3385, N93, N1550, N2410);
nand NAND4 (N3389, N3376, N2283, N49, N834);
nor NOR4 (N3390, N3359, N2002, N2611, N994);
not NOT1 (N3391, N3387);
nand NAND4 (N3392, N3372, N664, N1327, N1210);
nor NOR4 (N3393, N3389, N617, N529, N632);
not NOT1 (N3394, N3391);
buf BUF1 (N3395, N3381);
not NOT1 (N3396, N3382);
buf BUF1 (N3397, N3396);
nor NOR2 (N3398, N3397, N1069);
nor NOR3 (N3399, N3394, N2825, N2694);
not NOT1 (N3400, N3399);
buf BUF1 (N3401, N3386);
and AND2 (N3402, N3400, N1491);
buf BUF1 (N3403, N3395);
buf BUF1 (N3404, N3390);
nand NAND2 (N3405, N3404, N250);
and AND4 (N3406, N3402, N1761, N1883, N1477);
buf BUF1 (N3407, N3403);
xor XOR2 (N3408, N3398, N1674);
nand NAND4 (N3409, N3401, N2507, N2795, N1554);
not NOT1 (N3410, N3392);
or OR4 (N3411, N3408, N912, N2940, N443);
buf BUF1 (N3412, N3393);
and AND4 (N3413, N3383, N3142, N249, N1433);
buf BUF1 (N3414, N3407);
nor NOR4 (N3415, N3384, N160, N2306, N2079);
buf BUF1 (N3416, N3406);
xor XOR2 (N3417, N3415, N96);
xor XOR2 (N3418, N3417, N998);
nor NOR2 (N3419, N3413, N117);
or OR3 (N3420, N3411, N3395, N1102);
xor XOR2 (N3421, N3414, N13);
xor XOR2 (N3422, N3420, N1840);
buf BUF1 (N3423, N3388);
or OR3 (N3424, N3405, N2635, N76);
buf BUF1 (N3425, N3422);
nand NAND3 (N3426, N3421, N1137, N2172);
nor NOR2 (N3427, N3426, N2923);
nor NOR2 (N3428, N3425, N2504);
nor NOR3 (N3429, N3427, N1934, N2516);
or OR3 (N3430, N3418, N3429, N3102);
xor XOR2 (N3431, N991, N2260);
or OR3 (N3432, N3410, N2759, N1353);
or OR2 (N3433, N3409, N1225);
buf BUF1 (N3434, N3430);
not NOT1 (N3435, N3416);
nand NAND2 (N3436, N3412, N2233);
buf BUF1 (N3437, N3432);
xor XOR2 (N3438, N3437, N602);
xor XOR2 (N3439, N3428, N2821);
xor XOR2 (N3440, N3433, N3326);
nor NOR2 (N3441, N3434, N1411);
nor NOR2 (N3442, N3436, N315);
nand NAND4 (N3443, N3435, N1855, N2939, N324);
and AND4 (N3444, N3424, N2018, N2339, N2086);
buf BUF1 (N3445, N3440);
nor NOR2 (N3446, N3441, N2982);
buf BUF1 (N3447, N3423);
not NOT1 (N3448, N3445);
xor XOR2 (N3449, N3448, N2112);
buf BUF1 (N3450, N3438);
or OR3 (N3451, N3431, N3134, N1950);
nand NAND3 (N3452, N3439, N2051, N1273);
nand NAND3 (N3453, N3446, N1641, N2653);
and AND4 (N3454, N3453, N2985, N1568, N2449);
xor XOR2 (N3455, N3443, N662);
buf BUF1 (N3456, N3455);
and AND2 (N3457, N3456, N2651);
nand NAND3 (N3458, N3451, N84, N3369);
not NOT1 (N3459, N3450);
and AND2 (N3460, N3442, N2205);
and AND3 (N3461, N3454, N143, N2751);
xor XOR2 (N3462, N3447, N3346);
xor XOR2 (N3463, N3457, N2152);
not NOT1 (N3464, N3460);
nand NAND4 (N3465, N3449, N1252, N1600, N1557);
buf BUF1 (N3466, N3419);
xor XOR2 (N3467, N3461, N1445);
buf BUF1 (N3468, N3463);
nand NAND3 (N3469, N3452, N419, N710);
or OR3 (N3470, N3465, N2261, N2248);
and AND4 (N3471, N3468, N1913, N2406, N178);
and AND3 (N3472, N3469, N2386, N2400);
not NOT1 (N3473, N3462);
not NOT1 (N3474, N3444);
xor XOR2 (N3475, N3464, N2744);
nor NOR4 (N3476, N3471, N2768, N2603, N562);
or OR4 (N3477, N3473, N911, N733, N1510);
buf BUF1 (N3478, N3472);
nor NOR3 (N3479, N3477, N94, N848);
nor NOR2 (N3480, N3458, N895);
nand NAND2 (N3481, N3476, N491);
xor XOR2 (N3482, N3470, N548);
xor XOR2 (N3483, N3474, N1897);
buf BUF1 (N3484, N3483);
nor NOR2 (N3485, N3482, N3235);
nor NOR2 (N3486, N3480, N1011);
xor XOR2 (N3487, N3475, N1024);
buf BUF1 (N3488, N3459);
xor XOR2 (N3489, N3467, N1944);
or OR3 (N3490, N3489, N1439, N2968);
not NOT1 (N3491, N3487);
or OR4 (N3492, N3479, N2136, N2716, N3111);
nor NOR2 (N3493, N3466, N3006);
not NOT1 (N3494, N3490);
buf BUF1 (N3495, N3493);
xor XOR2 (N3496, N3495, N1575);
or OR2 (N3497, N3486, N301);
buf BUF1 (N3498, N3484);
buf BUF1 (N3499, N3492);
and AND4 (N3500, N3494, N921, N3154, N3469);
nand NAND4 (N3501, N3499, N1822, N180, N2775);
or OR4 (N3502, N3481, N1345, N804, N2396);
nand NAND3 (N3503, N3500, N2866, N680);
or OR4 (N3504, N3501, N1184, N686, N3348);
or OR3 (N3505, N3496, N1563, N3333);
or OR2 (N3506, N3498, N3190);
and AND4 (N3507, N3497, N2268, N722, N661);
nand NAND3 (N3508, N3485, N730, N1818);
nor NOR3 (N3509, N3506, N83, N1668);
buf BUF1 (N3510, N3478);
buf BUF1 (N3511, N3491);
and AND2 (N3512, N3488, N3272);
and AND3 (N3513, N3504, N2480, N2191);
or OR4 (N3514, N3511, N2588, N2763, N3288);
xor XOR2 (N3515, N3510, N561);
or OR2 (N3516, N3505, N575);
buf BUF1 (N3517, N3509);
or OR2 (N3518, N3515, N2015);
buf BUF1 (N3519, N3512);
nor NOR4 (N3520, N3513, N2449, N2652, N851);
nand NAND2 (N3521, N3507, N871);
xor XOR2 (N3522, N3518, N1676);
or OR2 (N3523, N3521, N3157);
and AND4 (N3524, N3520, N2929, N1173, N3258);
buf BUF1 (N3525, N3522);
or OR2 (N3526, N3514, N3317);
buf BUF1 (N3527, N3523);
and AND3 (N3528, N3517, N3290, N2500);
nand NAND4 (N3529, N3526, N2437, N214, N2853);
not NOT1 (N3530, N3519);
buf BUF1 (N3531, N3528);
and AND3 (N3532, N3503, N1066, N750);
or OR4 (N3533, N3525, N1360, N3391, N3222);
or OR4 (N3534, N3530, N1232, N3512, N1286);
and AND2 (N3535, N3516, N691);
or OR3 (N3536, N3535, N2948, N1731);
and AND3 (N3537, N3531, N2567, N1804);
and AND4 (N3538, N3502, N563, N2037, N908);
nand NAND3 (N3539, N3532, N821, N798);
not NOT1 (N3540, N3508);
or OR2 (N3541, N3536, N953);
nor NOR4 (N3542, N3537, N1077, N3131, N1523);
not NOT1 (N3543, N3527);
xor XOR2 (N3544, N3539, N1023);
nor NOR3 (N3545, N3543, N1484, N3307);
xor XOR2 (N3546, N3538, N1895);
not NOT1 (N3547, N3534);
and AND3 (N3548, N3544, N3384, N1588);
and AND4 (N3549, N3546, N350, N2362, N1887);
or OR2 (N3550, N3549, N114);
not NOT1 (N3551, N3540);
buf BUF1 (N3552, N3533);
not NOT1 (N3553, N3552);
or OR3 (N3554, N3524, N2417, N573);
nand NAND3 (N3555, N3545, N3511, N1915);
buf BUF1 (N3556, N3555);
and AND3 (N3557, N3529, N880, N69);
nand NAND3 (N3558, N3551, N1399, N607);
and AND3 (N3559, N3547, N3191, N3515);
buf BUF1 (N3560, N3553);
nand NAND2 (N3561, N3556, N1428);
not NOT1 (N3562, N3548);
xor XOR2 (N3563, N3558, N864);
nand NAND4 (N3564, N3562, N552, N708, N162);
and AND2 (N3565, N3550, N1715);
and AND4 (N3566, N3542, N3473, N2386, N1740);
and AND2 (N3567, N3561, N2792);
and AND2 (N3568, N3557, N3170);
buf BUF1 (N3569, N3554);
xor XOR2 (N3570, N3567, N1198);
buf BUF1 (N3571, N3560);
or OR2 (N3572, N3564, N3376);
and AND2 (N3573, N3569, N2463);
buf BUF1 (N3574, N3566);
and AND2 (N3575, N3571, N2864);
nor NOR2 (N3576, N3572, N2634);
and AND3 (N3577, N3570, N298, N2045);
nand NAND4 (N3578, N3573, N2374, N1146, N1354);
or OR3 (N3579, N3565, N1479, N3161);
nor NOR4 (N3580, N3563, N2055, N354, N3030);
and AND2 (N3581, N3580, N2248);
and AND2 (N3582, N3541, N77);
xor XOR2 (N3583, N3578, N732);
and AND4 (N3584, N3559, N924, N3465, N679);
nor NOR4 (N3585, N3584, N1008, N337, N3321);
nand NAND3 (N3586, N3583, N2718, N554);
not NOT1 (N3587, N3585);
xor XOR2 (N3588, N3568, N666);
not NOT1 (N3589, N3582);
xor XOR2 (N3590, N3586, N3090);
buf BUF1 (N3591, N3575);
buf BUF1 (N3592, N3590);
buf BUF1 (N3593, N3591);
xor XOR2 (N3594, N3574, N1871);
and AND2 (N3595, N3588, N2024);
nand NAND2 (N3596, N3577, N2508);
xor XOR2 (N3597, N3594, N2750);
nor NOR4 (N3598, N3596, N2948, N2731, N701);
or OR2 (N3599, N3593, N3276);
or OR2 (N3600, N3595, N1113);
buf BUF1 (N3601, N3599);
not NOT1 (N3602, N3587);
buf BUF1 (N3603, N3600);
xor XOR2 (N3604, N3576, N2609);
nor NOR2 (N3605, N3602, N2037);
nand NAND2 (N3606, N3592, N289);
buf BUF1 (N3607, N3604);
buf BUF1 (N3608, N3598);
or OR4 (N3609, N3603, N2933, N2083, N1152);
not NOT1 (N3610, N3589);
nand NAND3 (N3611, N3579, N1242, N1405);
nand NAND2 (N3612, N3607, N3440);
or OR4 (N3613, N3605, N2283, N399, N1198);
buf BUF1 (N3614, N3612);
not NOT1 (N3615, N3581);
not NOT1 (N3616, N3606);
nor NOR4 (N3617, N3616, N634, N2460, N929);
or OR2 (N3618, N3601, N2156);
nor NOR3 (N3619, N3597, N1913, N2218);
buf BUF1 (N3620, N3609);
nand NAND2 (N3621, N3617, N2333);
buf BUF1 (N3622, N3620);
or OR4 (N3623, N3615, N1003, N1738, N2752);
nand NAND2 (N3624, N3619, N335);
nand NAND4 (N3625, N3622, N58, N415, N3055);
nand NAND4 (N3626, N3624, N1675, N2886, N1874);
not NOT1 (N3627, N3614);
xor XOR2 (N3628, N3627, N1243);
or OR2 (N3629, N3628, N1859);
buf BUF1 (N3630, N3618);
nand NAND4 (N3631, N3625, N154, N2797, N2376);
and AND3 (N3632, N3629, N3071, N205);
not NOT1 (N3633, N3608);
or OR4 (N3634, N3633, N1867, N3257, N2674);
xor XOR2 (N3635, N3631, N2165);
buf BUF1 (N3636, N3611);
and AND3 (N3637, N3632, N2310, N503);
or OR4 (N3638, N3613, N1296, N226, N2675);
not NOT1 (N3639, N3636);
buf BUF1 (N3640, N3610);
buf BUF1 (N3641, N3639);
and AND2 (N3642, N3641, N633);
nor NOR3 (N3643, N3634, N755, N3560);
and AND4 (N3644, N3623, N2254, N1814, N977);
not NOT1 (N3645, N3642);
nor NOR2 (N3646, N3643, N2262);
nand NAND3 (N3647, N3640, N3539, N15);
or OR3 (N3648, N3630, N960, N3396);
buf BUF1 (N3649, N3647);
nor NOR2 (N3650, N3645, N2865);
nor NOR4 (N3651, N3626, N1381, N2512, N474);
not NOT1 (N3652, N3649);
or OR2 (N3653, N3644, N3536);
nor NOR2 (N3654, N3635, N2301);
buf BUF1 (N3655, N3651);
nand NAND3 (N3656, N3654, N1315, N3260);
nor NOR3 (N3657, N3646, N1403, N3134);
or OR4 (N3658, N3650, N1499, N1942, N2565);
xor XOR2 (N3659, N3648, N1354);
and AND3 (N3660, N3652, N815, N2939);
xor XOR2 (N3661, N3658, N1039);
or OR4 (N3662, N3621, N2389, N262, N1191);
not NOT1 (N3663, N3638);
and AND3 (N3664, N3656, N3151, N2508);
or OR2 (N3665, N3662, N83);
buf BUF1 (N3666, N3659);
and AND3 (N3667, N3664, N2560, N484);
xor XOR2 (N3668, N3655, N1908);
buf BUF1 (N3669, N3657);
xor XOR2 (N3670, N3668, N2809);
nand NAND2 (N3671, N3669, N3295);
nor NOR3 (N3672, N3665, N1133, N1921);
and AND3 (N3673, N3670, N2678, N1201);
and AND4 (N3674, N3660, N2591, N293, N1102);
buf BUF1 (N3675, N3653);
and AND3 (N3676, N3675, N2405, N730);
and AND4 (N3677, N3673, N1635, N612, N593);
xor XOR2 (N3678, N3671, N2636);
buf BUF1 (N3679, N3672);
and AND2 (N3680, N3667, N123);
or OR2 (N3681, N3637, N2388);
nand NAND4 (N3682, N3666, N3550, N1051, N2395);
buf BUF1 (N3683, N3679);
nor NOR3 (N3684, N3663, N328, N1661);
and AND2 (N3685, N3682, N848);
nand NAND2 (N3686, N3674, N1893);
buf BUF1 (N3687, N3684);
nand NAND2 (N3688, N3681, N824);
nand NAND2 (N3689, N3680, N1451);
buf BUF1 (N3690, N3686);
nand NAND4 (N3691, N3689, N3264, N1318, N2213);
nand NAND4 (N3692, N3691, N1949, N404, N108);
nor NOR4 (N3693, N3661, N402, N2955, N3685);
or OR4 (N3694, N3301, N1682, N456, N1437);
buf BUF1 (N3695, N3677);
buf BUF1 (N3696, N3692);
or OR2 (N3697, N3690, N2343);
nand NAND3 (N3698, N3693, N2570, N1365);
xor XOR2 (N3699, N3698, N716);
or OR2 (N3700, N3694, N1430);
nand NAND2 (N3701, N3688, N2695);
nor NOR3 (N3702, N3676, N1360, N1655);
nor NOR3 (N3703, N3696, N2164, N2565);
xor XOR2 (N3704, N3699, N1874);
or OR4 (N3705, N3702, N1090, N3071, N3526);
or OR3 (N3706, N3705, N1424, N3526);
not NOT1 (N3707, N3687);
and AND2 (N3708, N3704, N1629);
buf BUF1 (N3709, N3683);
buf BUF1 (N3710, N3709);
and AND2 (N3711, N3678, N3195);
not NOT1 (N3712, N3710);
xor XOR2 (N3713, N3711, N3212);
xor XOR2 (N3714, N3708, N1699);
or OR2 (N3715, N3706, N2165);
or OR2 (N3716, N3714, N1763);
buf BUF1 (N3717, N3707);
buf BUF1 (N3718, N3695);
nand NAND2 (N3719, N3713, N1956);
and AND4 (N3720, N3697, N3253, N3413, N1969);
xor XOR2 (N3721, N3718, N985);
nand NAND2 (N3722, N3716, N1568);
and AND3 (N3723, N3720, N2505, N3459);
nand NAND3 (N3724, N3721, N2469, N3349);
or OR4 (N3725, N3722, N2879, N1414, N3244);
buf BUF1 (N3726, N3719);
not NOT1 (N3727, N3726);
nor NOR4 (N3728, N3723, N80, N1283, N1688);
and AND2 (N3729, N3728, N2787);
not NOT1 (N3730, N3727);
or OR2 (N3731, N3725, N1277);
and AND4 (N3732, N3715, N19, N731, N5);
buf BUF1 (N3733, N3731);
buf BUF1 (N3734, N3730);
nor NOR4 (N3735, N3700, N2334, N2202, N1358);
nand NAND4 (N3736, N3701, N765, N2215, N2968);
or OR4 (N3737, N3703, N3339, N1531, N984);
nor NOR4 (N3738, N3737, N1312, N784, N2594);
not NOT1 (N3739, N3712);
not NOT1 (N3740, N3732);
nor NOR4 (N3741, N3734, N831, N687, N2641);
buf BUF1 (N3742, N3729);
nand NAND3 (N3743, N3735, N602, N2222);
and AND2 (N3744, N3741, N1328);
nor NOR2 (N3745, N3717, N1124);
not NOT1 (N3746, N3744);
nand NAND2 (N3747, N3733, N2154);
xor XOR2 (N3748, N3736, N1082);
or OR4 (N3749, N3747, N60, N120, N98);
xor XOR2 (N3750, N3746, N1196);
nor NOR2 (N3751, N3745, N2420);
not NOT1 (N3752, N3751);
xor XOR2 (N3753, N3738, N1091);
nor NOR4 (N3754, N3740, N283, N3456, N669);
buf BUF1 (N3755, N3752);
buf BUF1 (N3756, N3724);
and AND4 (N3757, N3754, N3516, N757, N3372);
and AND4 (N3758, N3739, N2476, N2641, N593);
or OR4 (N3759, N3749, N2739, N3323, N1897);
nor NOR4 (N3760, N3748, N1010, N3390, N87);
or OR3 (N3761, N3743, N1843, N402);
or OR4 (N3762, N3760, N1288, N1736, N1358);
nand NAND4 (N3763, N3753, N294, N409, N515);
or OR3 (N3764, N3755, N2905, N1713);
or OR3 (N3765, N3756, N2917, N53);
and AND4 (N3766, N3762, N469, N2187, N2739);
xor XOR2 (N3767, N3758, N598);
or OR4 (N3768, N3763, N2193, N2423, N2421);
not NOT1 (N3769, N3761);
xor XOR2 (N3770, N3750, N1086);
nor NOR3 (N3771, N3767, N1270, N1504);
or OR3 (N3772, N3768, N503, N3162);
not NOT1 (N3773, N3765);
and AND4 (N3774, N3766, N2420, N1777, N1776);
or OR2 (N3775, N3757, N3514);
buf BUF1 (N3776, N3764);
nor NOR2 (N3777, N3771, N989);
buf BUF1 (N3778, N3776);
not NOT1 (N3779, N3759);
nand NAND4 (N3780, N3773, N223, N446, N1342);
not NOT1 (N3781, N3772);
not NOT1 (N3782, N3780);
buf BUF1 (N3783, N3742);
not NOT1 (N3784, N3782);
buf BUF1 (N3785, N3777);
and AND3 (N3786, N3783, N3042, N2345);
not NOT1 (N3787, N3784);
not NOT1 (N3788, N3778);
nor NOR2 (N3789, N3786, N2822);
buf BUF1 (N3790, N3789);
xor XOR2 (N3791, N3775, N3659);
nand NAND4 (N3792, N3791, N1038, N3694, N868);
and AND2 (N3793, N3792, N1881);
xor XOR2 (N3794, N3790, N240);
nor NOR3 (N3795, N3769, N1441, N3009);
nand NAND3 (N3796, N3788, N1318, N1024);
xor XOR2 (N3797, N3795, N3249);
xor XOR2 (N3798, N3781, N424);
xor XOR2 (N3799, N3797, N2677);
xor XOR2 (N3800, N3785, N2684);
xor XOR2 (N3801, N3799, N1589);
and AND2 (N3802, N3794, N633);
not NOT1 (N3803, N3774);
not NOT1 (N3804, N3801);
buf BUF1 (N3805, N3798);
or OR3 (N3806, N3802, N1281, N998);
nor NOR3 (N3807, N3779, N2129, N169);
buf BUF1 (N3808, N3787);
buf BUF1 (N3809, N3800);
nand NAND3 (N3810, N3804, N1152, N170);
buf BUF1 (N3811, N3809);
nand NAND3 (N3812, N3770, N1938, N3283);
or OR2 (N3813, N3807, N3089);
not NOT1 (N3814, N3793);
and AND3 (N3815, N3805, N3288, N1325);
not NOT1 (N3816, N3813);
or OR2 (N3817, N3810, N627);
or OR2 (N3818, N3814, N1372);
xor XOR2 (N3819, N3818, N3780);
xor XOR2 (N3820, N3815, N1412);
xor XOR2 (N3821, N3811, N3607);
or OR2 (N3822, N3806, N985);
buf BUF1 (N3823, N3819);
nand NAND2 (N3824, N3812, N1459);
buf BUF1 (N3825, N3817);
buf BUF1 (N3826, N3816);
and AND3 (N3827, N3825, N279, N3064);
buf BUF1 (N3828, N3826);
or OR4 (N3829, N3827, N1150, N613, N2938);
xor XOR2 (N3830, N3803, N3589);
not NOT1 (N3831, N3796);
xor XOR2 (N3832, N3831, N1024);
and AND4 (N3833, N3823, N400, N2378, N3468);
nor NOR2 (N3834, N3828, N2182);
buf BUF1 (N3835, N3834);
buf BUF1 (N3836, N3833);
nand NAND2 (N3837, N3824, N3045);
or OR3 (N3838, N3820, N20, N1257);
not NOT1 (N3839, N3829);
not NOT1 (N3840, N3821);
buf BUF1 (N3841, N3832);
or OR3 (N3842, N3839, N2219, N2989);
nor NOR4 (N3843, N3808, N3762, N2579, N1319);
or OR2 (N3844, N3838, N2999);
or OR2 (N3845, N3844, N1617);
xor XOR2 (N3846, N3842, N1862);
nand NAND2 (N3847, N3846, N1319);
buf BUF1 (N3848, N3845);
and AND2 (N3849, N3822, N1494);
or OR2 (N3850, N3849, N1636);
buf BUF1 (N3851, N3836);
not NOT1 (N3852, N3850);
xor XOR2 (N3853, N3837, N2154);
buf BUF1 (N3854, N3843);
and AND3 (N3855, N3851, N973, N1540);
not NOT1 (N3856, N3855);
nand NAND2 (N3857, N3841, N2617);
xor XOR2 (N3858, N3848, N2330);
buf BUF1 (N3859, N3847);
or OR4 (N3860, N3858, N1309, N1705, N3373);
not NOT1 (N3861, N3859);
buf BUF1 (N3862, N3830);
not NOT1 (N3863, N3840);
xor XOR2 (N3864, N3853, N1186);
buf BUF1 (N3865, N3854);
or OR3 (N3866, N3861, N2358, N3466);
nor NOR2 (N3867, N3860, N217);
and AND2 (N3868, N3852, N2829);
buf BUF1 (N3869, N3867);
buf BUF1 (N3870, N3862);
nor NOR4 (N3871, N3864, N3669, N1167, N1646);
not NOT1 (N3872, N3869);
buf BUF1 (N3873, N3857);
nor NOR2 (N3874, N3866, N779);
xor XOR2 (N3875, N3865, N3557);
nand NAND4 (N3876, N3835, N631, N2236, N1696);
nor NOR4 (N3877, N3873, N3246, N3072, N791);
nor NOR2 (N3878, N3863, N3268);
xor XOR2 (N3879, N3868, N3218);
and AND3 (N3880, N3856, N190, N3655);
nor NOR4 (N3881, N3871, N2245, N1526, N3439);
nand NAND4 (N3882, N3870, N3122, N1681, N1466);
or OR2 (N3883, N3877, N3755);
nor NOR4 (N3884, N3876, N1449, N949, N864);
and AND3 (N3885, N3883, N1081, N3716);
nand NAND3 (N3886, N3880, N3843, N3324);
nor NOR3 (N3887, N3878, N3864, N1666);
or OR2 (N3888, N3884, N3186);
or OR2 (N3889, N3887, N1752);
not NOT1 (N3890, N3874);
nor NOR3 (N3891, N3872, N2741, N1441);
xor XOR2 (N3892, N3881, N2200);
xor XOR2 (N3893, N3885, N2157);
or OR3 (N3894, N3890, N2531, N1067);
xor XOR2 (N3895, N3891, N3308);
and AND4 (N3896, N3892, N2605, N2579, N3003);
and AND3 (N3897, N3879, N36, N3321);
nor NOR2 (N3898, N3882, N48);
and AND2 (N3899, N3898, N1005);
not NOT1 (N3900, N3888);
and AND2 (N3901, N3893, N2876);
buf BUF1 (N3902, N3896);
xor XOR2 (N3903, N3897, N1897);
buf BUF1 (N3904, N3903);
xor XOR2 (N3905, N3875, N934);
or OR2 (N3906, N3894, N3059);
buf BUF1 (N3907, N3902);
not NOT1 (N3908, N3889);
not NOT1 (N3909, N3908);
xor XOR2 (N3910, N3905, N1830);
not NOT1 (N3911, N3906);
nor NOR2 (N3912, N3886, N578);
nor NOR4 (N3913, N3904, N1047, N2921, N440);
or OR4 (N3914, N3911, N1994, N640, N170);
and AND4 (N3915, N3914, N264, N1452, N825);
buf BUF1 (N3916, N3910);
nor NOR3 (N3917, N3907, N3367, N2760);
or OR4 (N3918, N3909, N989, N642, N770);
not NOT1 (N3919, N3916);
or OR4 (N3920, N3901, N1753, N2758, N1945);
or OR4 (N3921, N3920, N2375, N327, N2429);
buf BUF1 (N3922, N3918);
not NOT1 (N3923, N3917);
nor NOR3 (N3924, N3922, N1487, N1387);
nor NOR3 (N3925, N3899, N2596, N658);
not NOT1 (N3926, N3921);
and AND2 (N3927, N3912, N2175);
or OR4 (N3928, N3926, N1831, N1839, N2505);
not NOT1 (N3929, N3924);
buf BUF1 (N3930, N3915);
buf BUF1 (N3931, N3925);
nand NAND4 (N3932, N3928, N3154, N2686, N3665);
nor NOR4 (N3933, N3931, N2213, N3050, N3171);
buf BUF1 (N3934, N3913);
xor XOR2 (N3935, N3923, N1667);
and AND4 (N3936, N3927, N2627, N2284, N3367);
buf BUF1 (N3937, N3932);
xor XOR2 (N3938, N3930, N909);
xor XOR2 (N3939, N3936, N1127);
and AND2 (N3940, N3938, N34);
nor NOR2 (N3941, N3940, N1743);
nand NAND4 (N3942, N3919, N1842, N1499, N2723);
buf BUF1 (N3943, N3895);
nand NAND4 (N3944, N3933, N3374, N691, N3799);
nor NOR2 (N3945, N3944, N885);
nand NAND4 (N3946, N3941, N3296, N2926, N2055);
or OR2 (N3947, N3934, N2885);
and AND3 (N3948, N3946, N220, N1162);
nand NAND4 (N3949, N3948, N3716, N423, N3051);
buf BUF1 (N3950, N3935);
or OR3 (N3951, N3900, N800, N63);
and AND4 (N3952, N3949, N870, N3604, N1809);
and AND4 (N3953, N3947, N1513, N2769, N345);
nand NAND2 (N3954, N3929, N2739);
not NOT1 (N3955, N3943);
not NOT1 (N3956, N3952);
buf BUF1 (N3957, N3956);
xor XOR2 (N3958, N3942, N615);
and AND2 (N3959, N3955, N202);
not NOT1 (N3960, N3953);
or OR3 (N3961, N3937, N3100, N3519);
or OR3 (N3962, N3951, N3896, N3755);
nand NAND3 (N3963, N3939, N2766, N3263);
buf BUF1 (N3964, N3950);
nand NAND4 (N3965, N3962, N2806, N315, N1285);
or OR2 (N3966, N3954, N730);
nand NAND2 (N3967, N3959, N3144);
buf BUF1 (N3968, N3965);
nor NOR2 (N3969, N3966, N3762);
and AND2 (N3970, N3961, N2665);
nor NOR2 (N3971, N3957, N3774);
or OR2 (N3972, N3945, N2872);
or OR3 (N3973, N3968, N2336, N3780);
and AND2 (N3974, N3967, N460);
xor XOR2 (N3975, N3963, N1811);
not NOT1 (N3976, N3975);
nand NAND2 (N3977, N3976, N3185);
and AND2 (N3978, N3972, N300);
and AND2 (N3979, N3964, N1328);
and AND3 (N3980, N3970, N22, N1663);
or OR2 (N3981, N3978, N2345);
and AND2 (N3982, N3958, N3454);
nor NOR4 (N3983, N3979, N3861, N3702, N354);
not NOT1 (N3984, N3974);
and AND2 (N3985, N3982, N1174);
nand NAND4 (N3986, N3971, N1687, N2305, N3529);
and AND2 (N3987, N3985, N3305);
nor NOR3 (N3988, N3973, N2463, N276);
xor XOR2 (N3989, N3977, N3041);
buf BUF1 (N3990, N3980);
nand NAND3 (N3991, N3983, N1285, N3500);
xor XOR2 (N3992, N3960, N3427);
xor XOR2 (N3993, N3990, N3027);
buf BUF1 (N3994, N3991);
and AND4 (N3995, N3992, N189, N3748, N114);
nand NAND3 (N3996, N3986, N3554, N1137);
buf BUF1 (N3997, N3984);
or OR2 (N3998, N3997, N1230);
and AND3 (N3999, N3993, N2895, N300);
nand NAND2 (N4000, N3994, N2774);
buf BUF1 (N4001, N3969);
or OR4 (N4002, N3999, N2236, N2868, N2370);
or OR3 (N4003, N4000, N634, N801);
xor XOR2 (N4004, N3987, N2340);
xor XOR2 (N4005, N3989, N278);
nand NAND2 (N4006, N3996, N4005);
buf BUF1 (N4007, N3608);
buf BUF1 (N4008, N4007);
or OR2 (N4009, N4001, N1501);
and AND2 (N4010, N4006, N804);
xor XOR2 (N4011, N4004, N1105);
or OR2 (N4012, N4010, N332);
nor NOR2 (N4013, N3988, N2603);
buf BUF1 (N4014, N4002);
or OR2 (N4015, N4012, N610);
or OR2 (N4016, N4014, N1628);
buf BUF1 (N4017, N3981);
nor NOR3 (N4018, N4017, N385, N3406);
not NOT1 (N4019, N3995);
xor XOR2 (N4020, N4008, N1462);
not NOT1 (N4021, N4018);
nor NOR4 (N4022, N4020, N1952, N1358, N1157);
nand NAND2 (N4023, N4003, N1837);
xor XOR2 (N4024, N4019, N3419);
or OR4 (N4025, N4024, N466, N1232, N2845);
nor NOR4 (N4026, N4016, N1347, N1896, N3137);
xor XOR2 (N4027, N4013, N2841);
nand NAND2 (N4028, N4021, N2415);
xor XOR2 (N4029, N4025, N286);
xor XOR2 (N4030, N4027, N767);
and AND3 (N4031, N4015, N365, N3626);
and AND4 (N4032, N4031, N3179, N577, N1796);
xor XOR2 (N4033, N4026, N1969);
xor XOR2 (N4034, N4029, N119);
nor NOR4 (N4035, N3998, N3402, N1510, N2729);
and AND3 (N4036, N4033, N2081, N1781);
not NOT1 (N4037, N4022);
xor XOR2 (N4038, N4037, N2663);
nor NOR2 (N4039, N4023, N621);
buf BUF1 (N4040, N4011);
buf BUF1 (N4041, N4038);
xor XOR2 (N4042, N4035, N2706);
and AND4 (N4043, N4032, N3121, N1199, N3828);
and AND2 (N4044, N4034, N3595);
buf BUF1 (N4045, N4028);
nor NOR4 (N4046, N4009, N1493, N3580, N2245);
or OR3 (N4047, N4040, N2265, N3266);
nand NAND2 (N4048, N4036, N3810);
and AND2 (N4049, N4041, N298);
buf BUF1 (N4050, N4043);
nor NOR2 (N4051, N4048, N2439);
and AND4 (N4052, N4050, N3344, N1907, N288);
xor XOR2 (N4053, N4030, N2451);
xor XOR2 (N4054, N4039, N3064);
and AND4 (N4055, N4042, N939, N3229, N1174);
or OR3 (N4056, N4047, N261, N1950);
nor NOR2 (N4057, N4051, N1498);
xor XOR2 (N4058, N4056, N165);
nand NAND4 (N4059, N4053, N2959, N3850, N1027);
nor NOR4 (N4060, N4049, N3606, N908, N3441);
or OR4 (N4061, N4045, N1365, N1587, N3573);
nand NAND2 (N4062, N4060, N1823);
nor NOR4 (N4063, N4054, N3466, N622, N222);
or OR2 (N4064, N4044, N453);
xor XOR2 (N4065, N4052, N511);
or OR4 (N4066, N4062, N3973, N3279, N3375);
not NOT1 (N4067, N4066);
nand NAND4 (N4068, N4067, N1731, N2507, N2023);
or OR2 (N4069, N4064, N1477);
nand NAND4 (N4070, N4065, N1196, N2616, N914);
not NOT1 (N4071, N4061);
buf BUF1 (N4072, N4055);
nand NAND2 (N4073, N4063, N1097);
nor NOR3 (N4074, N4059, N2522, N2893);
or OR4 (N4075, N4072, N1594, N958, N175);
and AND2 (N4076, N4068, N3248);
and AND3 (N4077, N4075, N2664, N1799);
nand NAND4 (N4078, N4076, N1490, N465, N2601);
xor XOR2 (N4079, N4069, N752);
and AND4 (N4080, N4057, N2839, N2863, N1587);
not NOT1 (N4081, N4077);
nor NOR3 (N4082, N4058, N2714, N751);
not NOT1 (N4083, N4046);
or OR2 (N4084, N4081, N548);
not NOT1 (N4085, N4070);
nor NOR3 (N4086, N4082, N3412, N1304);
xor XOR2 (N4087, N4078, N2000);
nand NAND3 (N4088, N4079, N1714, N972);
buf BUF1 (N4089, N4085);
xor XOR2 (N4090, N4088, N3993);
buf BUF1 (N4091, N4071);
and AND3 (N4092, N4089, N1386, N1112);
nor NOR2 (N4093, N4074, N913);
nor NOR2 (N4094, N4083, N148);
nand NAND3 (N4095, N4084, N3598, N3401);
nand NAND3 (N4096, N4086, N3260, N40);
or OR4 (N4097, N4087, N3543, N991, N3194);
or OR3 (N4098, N4090, N476, N1887);
nand NAND4 (N4099, N4098, N1966, N866, N1572);
nand NAND2 (N4100, N4096, N189);
not NOT1 (N4101, N4092);
and AND2 (N4102, N4093, N2359);
not NOT1 (N4103, N4101);
or OR3 (N4104, N4080, N2106, N3827);
not NOT1 (N4105, N4104);
and AND2 (N4106, N4100, N920);
xor XOR2 (N4107, N4102, N2230);
buf BUF1 (N4108, N4103);
nor NOR3 (N4109, N4108, N1880, N1011);
and AND4 (N4110, N4073, N2993, N1093, N3638);
and AND4 (N4111, N4106, N949, N2842, N1326);
xor XOR2 (N4112, N4094, N1711);
nor NOR2 (N4113, N4111, N1746);
and AND4 (N4114, N4112, N3819, N2066, N242);
nor NOR3 (N4115, N4095, N1727, N394);
or OR3 (N4116, N4091, N3025, N3297);
nand NAND3 (N4117, N4110, N2173, N3146);
not NOT1 (N4118, N4097);
and AND3 (N4119, N4109, N3727, N2997);
not NOT1 (N4120, N4113);
nand NAND2 (N4121, N4119, N2920);
buf BUF1 (N4122, N4120);
not NOT1 (N4123, N4122);
xor XOR2 (N4124, N4121, N1271);
xor XOR2 (N4125, N4107, N1491);
not NOT1 (N4126, N4123);
nand NAND3 (N4127, N4114, N3963, N295);
nor NOR3 (N4128, N4124, N3045, N2768);
buf BUF1 (N4129, N4128);
nor NOR4 (N4130, N4115, N1776, N2853, N1357);
buf BUF1 (N4131, N4105);
not NOT1 (N4132, N4116);
and AND2 (N4133, N4099, N3516);
buf BUF1 (N4134, N4118);
not NOT1 (N4135, N4132);
buf BUF1 (N4136, N4129);
nor NOR3 (N4137, N4131, N1931, N3249);
nor NOR2 (N4138, N4135, N1769);
or OR4 (N4139, N4126, N2102, N2416, N891);
xor XOR2 (N4140, N4117, N3105);
and AND4 (N4141, N4125, N2127, N394, N416);
nand NAND2 (N4142, N4137, N2970);
or OR3 (N4143, N4142, N1770, N1505);
nand NAND2 (N4144, N4130, N3784);
and AND4 (N4145, N4139, N3632, N3791, N1378);
or OR2 (N4146, N4141, N1462);
nand NAND2 (N4147, N4140, N13);
nand NAND3 (N4148, N4133, N3340, N1167);
nor NOR3 (N4149, N4144, N3353, N2782);
buf BUF1 (N4150, N4149);
buf BUF1 (N4151, N4148);
nand NAND2 (N4152, N4127, N2427);
or OR4 (N4153, N4136, N3300, N1112, N3217);
xor XOR2 (N4154, N4143, N2449);
nor NOR2 (N4155, N4151, N2605);
xor XOR2 (N4156, N4146, N4129);
nor NOR4 (N4157, N4154, N2740, N1433, N1321);
xor XOR2 (N4158, N4156, N105);
nor NOR4 (N4159, N4147, N1679, N1351, N380);
nand NAND2 (N4160, N4153, N2180);
not NOT1 (N4161, N4134);
and AND2 (N4162, N4158, N1825);
nand NAND3 (N4163, N4152, N4092, N179);
or OR4 (N4164, N4160, N4032, N3424, N8);
nor NOR2 (N4165, N4164, N1589);
nand NAND3 (N4166, N4155, N4102, N131);
nor NOR3 (N4167, N4166, N555, N235);
buf BUF1 (N4168, N4162);
xor XOR2 (N4169, N4163, N46);
xor XOR2 (N4170, N4138, N1659);
buf BUF1 (N4171, N4157);
nand NAND3 (N4172, N4169, N3854, N2772);
nor NOR4 (N4173, N4167, N1958, N1338, N1937);
and AND4 (N4174, N4170, N1488, N3670, N4045);
or OR2 (N4175, N4145, N2426);
xor XOR2 (N4176, N4168, N2255);
or OR2 (N4177, N4175, N3500);
and AND4 (N4178, N4176, N1715, N3940, N806);
nor NOR2 (N4179, N4172, N3197);
nor NOR3 (N4180, N4161, N1558, N1090);
or OR3 (N4181, N4179, N2586, N3334);
not NOT1 (N4182, N4171);
or OR3 (N4183, N4165, N837, N1084);
not NOT1 (N4184, N4150);
not NOT1 (N4185, N4177);
nand NAND3 (N4186, N4180, N3073, N1559);
buf BUF1 (N4187, N4174);
or OR3 (N4188, N4159, N1441, N3191);
nand NAND3 (N4189, N4185, N65, N1665);
nand NAND2 (N4190, N4182, N767);
buf BUF1 (N4191, N4187);
nand NAND4 (N4192, N4188, N1885, N2449, N3747);
xor XOR2 (N4193, N4190, N2455);
nor NOR4 (N4194, N4191, N1777, N3287, N214);
not NOT1 (N4195, N4178);
nand NAND3 (N4196, N4186, N1241, N40);
nor NOR3 (N4197, N4196, N71, N1637);
and AND2 (N4198, N4183, N1641);
nand NAND2 (N4199, N4189, N2493);
xor XOR2 (N4200, N4181, N1409);
xor XOR2 (N4201, N4198, N3138);
xor XOR2 (N4202, N4192, N3315);
not NOT1 (N4203, N4201);
or OR2 (N4204, N4199, N3139);
nor NOR4 (N4205, N4193, N1500, N3133, N1527);
xor XOR2 (N4206, N4205, N351);
nor NOR2 (N4207, N4173, N1074);
and AND3 (N4208, N4204, N1180, N404);
nor NOR2 (N4209, N4202, N3702);
buf BUF1 (N4210, N4197);
xor XOR2 (N4211, N4203, N851);
buf BUF1 (N4212, N4207);
not NOT1 (N4213, N4206);
nor NOR3 (N4214, N4210, N2237, N1740);
or OR4 (N4215, N4200, N2610, N601, N2047);
not NOT1 (N4216, N4208);
and AND4 (N4217, N4212, N225, N884, N3383);
not NOT1 (N4218, N4215);
xor XOR2 (N4219, N4218, N86);
or OR2 (N4220, N4213, N643);
xor XOR2 (N4221, N4220, N618);
buf BUF1 (N4222, N4195);
and AND4 (N4223, N4194, N1673, N205, N3603);
xor XOR2 (N4224, N4184, N989);
xor XOR2 (N4225, N4221, N1255);
or OR2 (N4226, N4224, N2202);
nand NAND4 (N4227, N4211, N3096, N1334, N2341);
xor XOR2 (N4228, N4216, N3540);
nor NOR2 (N4229, N4225, N3138);
and AND3 (N4230, N4214, N3467, N1978);
not NOT1 (N4231, N4226);
buf BUF1 (N4232, N4228);
buf BUF1 (N4233, N4229);
xor XOR2 (N4234, N4222, N3022);
buf BUF1 (N4235, N4219);
or OR2 (N4236, N4233, N3813);
nor NOR4 (N4237, N4232, N2833, N790, N3518);
or OR3 (N4238, N4234, N1168, N2295);
nand NAND2 (N4239, N4231, N3139);
nand NAND2 (N4240, N4230, N3670);
xor XOR2 (N4241, N4239, N263);
and AND2 (N4242, N4209, N2802);
or OR3 (N4243, N4240, N724, N3972);
and AND2 (N4244, N4243, N2868);
nand NAND4 (N4245, N4242, N2104, N1145, N3613);
or OR2 (N4246, N4217, N3932);
and AND2 (N4247, N4223, N467);
xor XOR2 (N4248, N4247, N222);
or OR3 (N4249, N4245, N2321, N3802);
and AND2 (N4250, N4238, N1048);
and AND2 (N4251, N4250, N230);
nand NAND2 (N4252, N4235, N196);
or OR4 (N4253, N4252, N1932, N1474, N2635);
buf BUF1 (N4254, N4236);
nor NOR2 (N4255, N4227, N2427);
and AND3 (N4256, N4251, N2623, N3934);
nand NAND3 (N4257, N4246, N3559, N2857);
or OR3 (N4258, N4237, N797, N3602);
and AND2 (N4259, N4249, N2873);
xor XOR2 (N4260, N4244, N2631);
xor XOR2 (N4261, N4258, N2899);
xor XOR2 (N4262, N4241, N4120);
buf BUF1 (N4263, N4261);
or OR2 (N4264, N4262, N1926);
not NOT1 (N4265, N4255);
buf BUF1 (N4266, N4248);
or OR3 (N4267, N4259, N874, N549);
buf BUF1 (N4268, N4263);
xor XOR2 (N4269, N4260, N673);
xor XOR2 (N4270, N4268, N309);
or OR2 (N4271, N4270, N4061);
buf BUF1 (N4272, N4256);
xor XOR2 (N4273, N4253, N27);
xor XOR2 (N4274, N4254, N3266);
not NOT1 (N4275, N4267);
not NOT1 (N4276, N4264);
nand NAND3 (N4277, N4274, N3565, N4002);
or OR2 (N4278, N4265, N3994);
buf BUF1 (N4279, N4275);
not NOT1 (N4280, N4272);
and AND2 (N4281, N4277, N2808);
or OR4 (N4282, N4269, N4218, N3153, N395);
and AND3 (N4283, N4281, N1184, N1935);
nand NAND2 (N4284, N4282, N559);
and AND2 (N4285, N4271, N2375);
or OR2 (N4286, N4284, N231);
nand NAND2 (N4287, N4286, N277);
not NOT1 (N4288, N4273);
nor NOR2 (N4289, N4288, N2881);
not NOT1 (N4290, N4285);
nor NOR4 (N4291, N4278, N2178, N356, N3404);
buf BUF1 (N4292, N4291);
buf BUF1 (N4293, N4280);
nor NOR2 (N4294, N4279, N2836);
nor NOR4 (N4295, N4293, N1965, N4128, N2775);
buf BUF1 (N4296, N4295);
nor NOR2 (N4297, N4287, N169);
buf BUF1 (N4298, N4257);
or OR3 (N4299, N4290, N258, N417);
or OR2 (N4300, N4299, N397);
buf BUF1 (N4301, N4294);
xor XOR2 (N4302, N4266, N3193);
nor NOR4 (N4303, N4292, N3751, N3142, N1881);
nor NOR3 (N4304, N4296, N1000, N747);
xor XOR2 (N4305, N4303, N323);
nand NAND3 (N4306, N4304, N2221, N43);
or OR4 (N4307, N4276, N2913, N3914, N1410);
or OR3 (N4308, N4300, N2368, N3171);
nor NOR4 (N4309, N4306, N1085, N2537, N1685);
or OR4 (N4310, N4297, N1020, N1916, N2577);
nor NOR2 (N4311, N4301, N2160);
nand NAND4 (N4312, N4283, N2578, N744, N1297);
nor NOR3 (N4313, N4289, N2558, N3939);
xor XOR2 (N4314, N4305, N3944);
buf BUF1 (N4315, N4311);
xor XOR2 (N4316, N4310, N3733);
nand NAND2 (N4317, N4316, N2568);
xor XOR2 (N4318, N4309, N2861);
xor XOR2 (N4319, N4298, N1916);
xor XOR2 (N4320, N4319, N561);
nand NAND4 (N4321, N4314, N4267, N3691, N1469);
nor NOR4 (N4322, N4320, N173, N1061, N2427);
xor XOR2 (N4323, N4322, N1493);
buf BUF1 (N4324, N4315);
not NOT1 (N4325, N4308);
xor XOR2 (N4326, N4312, N1713);
nand NAND2 (N4327, N4313, N3316);
or OR4 (N4328, N4317, N402, N2801, N2559);
nand NAND2 (N4329, N4327, N2164);
nor NOR2 (N4330, N4328, N163);
nor NOR3 (N4331, N4318, N2540, N3201);
nand NAND2 (N4332, N4324, N1960);
or OR4 (N4333, N4321, N289, N2911, N4228);
buf BUF1 (N4334, N4332);
not NOT1 (N4335, N4307);
and AND2 (N4336, N4325, N3032);
buf BUF1 (N4337, N4333);
buf BUF1 (N4338, N4337);
and AND3 (N4339, N4323, N3689, N3954);
buf BUF1 (N4340, N4339);
buf BUF1 (N4341, N4338);
nor NOR3 (N4342, N4340, N1938, N531);
or OR2 (N4343, N4329, N474);
and AND3 (N4344, N4342, N2386, N1146);
and AND3 (N4345, N4302, N1577, N159);
xor XOR2 (N4346, N4335, N2541);
not NOT1 (N4347, N4334);
not NOT1 (N4348, N4341);
xor XOR2 (N4349, N4331, N3489);
nor NOR4 (N4350, N4326, N1924, N3003, N800);
and AND2 (N4351, N4346, N4019);
buf BUF1 (N4352, N4343);
and AND3 (N4353, N4350, N3089, N3509);
nor NOR2 (N4354, N4330, N2124);
or OR2 (N4355, N4347, N1602);
or OR2 (N4356, N4354, N3083);
or OR2 (N4357, N4349, N3950);
buf BUF1 (N4358, N4348);
or OR2 (N4359, N4336, N895);
or OR4 (N4360, N4358, N3585, N2168, N581);
xor XOR2 (N4361, N4352, N682);
nor NOR3 (N4362, N4360, N487, N1702);
not NOT1 (N4363, N4362);
not NOT1 (N4364, N4357);
nor NOR2 (N4365, N4361, N3768);
nand NAND3 (N4366, N4345, N2750, N1270);
and AND3 (N4367, N4355, N2146, N2644);
nand NAND4 (N4368, N4365, N73, N581, N1310);
not NOT1 (N4369, N4359);
xor XOR2 (N4370, N4367, N140);
nor NOR2 (N4371, N4344, N2533);
not NOT1 (N4372, N4353);
not NOT1 (N4373, N4370);
nor NOR3 (N4374, N4366, N879, N2233);
xor XOR2 (N4375, N4372, N1835);
not NOT1 (N4376, N4371);
not NOT1 (N4377, N4376);
nor NOR4 (N4378, N4373, N4026, N3082, N4346);
nor NOR4 (N4379, N4377, N3796, N534, N2481);
not NOT1 (N4380, N4363);
buf BUF1 (N4381, N4374);
and AND4 (N4382, N4369, N1110, N454, N2860);
xor XOR2 (N4383, N4356, N2573);
nor NOR2 (N4384, N4381, N1923);
nor NOR4 (N4385, N4351, N4347, N580, N4215);
buf BUF1 (N4386, N4382);
or OR3 (N4387, N4364, N286, N3308);
nor NOR2 (N4388, N4385, N4028);
or OR2 (N4389, N4378, N1920);
xor XOR2 (N4390, N4386, N64);
buf BUF1 (N4391, N4383);
not NOT1 (N4392, N4391);
buf BUF1 (N4393, N4390);
buf BUF1 (N4394, N4368);
or OR4 (N4395, N4387, N2314, N3218, N621);
not NOT1 (N4396, N4380);
not NOT1 (N4397, N4393);
buf BUF1 (N4398, N4375);
and AND4 (N4399, N4397, N2221, N4220, N1799);
buf BUF1 (N4400, N4395);
or OR3 (N4401, N4388, N189, N1742);
not NOT1 (N4402, N4401);
and AND4 (N4403, N4394, N65, N2822, N4282);
or OR3 (N4404, N4403, N1351, N1029);
or OR3 (N4405, N4392, N1355, N2222);
buf BUF1 (N4406, N4384);
not NOT1 (N4407, N4399);
xor XOR2 (N4408, N4404, N1622);
and AND3 (N4409, N4405, N41, N591);
and AND2 (N4410, N4398, N429);
or OR3 (N4411, N4410, N470, N141);
nor NOR3 (N4412, N4409, N2307, N3487);
buf BUF1 (N4413, N4402);
or OR3 (N4414, N4406, N1279, N3241);
or OR4 (N4415, N4407, N2727, N2900, N989);
nand NAND4 (N4416, N4412, N1476, N309, N2437);
or OR4 (N4417, N4414, N2109, N2660, N2551);
and AND4 (N4418, N4379, N3897, N3907, N2908);
or OR3 (N4419, N4400, N3442, N1830);
xor XOR2 (N4420, N4408, N377);
or OR4 (N4421, N4415, N3963, N2508, N2064);
or OR3 (N4422, N4389, N4295, N4245);
and AND2 (N4423, N4418, N407);
and AND2 (N4424, N4396, N2718);
buf BUF1 (N4425, N4411);
xor XOR2 (N4426, N4422, N1508);
nand NAND2 (N4427, N4421, N2870);
and AND4 (N4428, N4425, N476, N3406, N4213);
or OR2 (N4429, N4417, N543);
not NOT1 (N4430, N4420);
not NOT1 (N4431, N4427);
not NOT1 (N4432, N4419);
and AND2 (N4433, N4428, N1859);
or OR2 (N4434, N4431, N3246);
not NOT1 (N4435, N4430);
or OR2 (N4436, N4433, N3407);
nor NOR2 (N4437, N4429, N840);
not NOT1 (N4438, N4432);
nand NAND2 (N4439, N4424, N1732);
and AND2 (N4440, N4423, N1357);
nand NAND2 (N4441, N4426, N2993);
nand NAND3 (N4442, N4413, N2710, N1614);
buf BUF1 (N4443, N4439);
not NOT1 (N4444, N4434);
nand NAND4 (N4445, N4416, N1766, N1089, N241);
buf BUF1 (N4446, N4443);
not NOT1 (N4447, N4442);
nor NOR4 (N4448, N4447, N1756, N3803, N146);
not NOT1 (N4449, N4440);
not NOT1 (N4450, N4449);
not NOT1 (N4451, N4445);
buf BUF1 (N4452, N4444);
buf BUF1 (N4453, N4446);
or OR2 (N4454, N4448, N1136);
or OR2 (N4455, N4437, N522);
and AND4 (N4456, N4441, N3291, N1209, N1607);
nor NOR4 (N4457, N4455, N916, N3395, N2014);
nor NOR4 (N4458, N4435, N1862, N2415, N4300);
buf BUF1 (N4459, N4453);
and AND2 (N4460, N4438, N1672);
nor NOR2 (N4461, N4456, N2945);
nand NAND2 (N4462, N4460, N319);
not NOT1 (N4463, N4454);
nand NAND2 (N4464, N4463, N546);
nand NAND4 (N4465, N4459, N2072, N3114, N2397);
xor XOR2 (N4466, N4450, N1256);
xor XOR2 (N4467, N4452, N4063);
not NOT1 (N4468, N4458);
and AND4 (N4469, N4464, N2769, N1488, N2824);
xor XOR2 (N4470, N4461, N3125);
buf BUF1 (N4471, N4462);
not NOT1 (N4472, N4457);
nor NOR3 (N4473, N4469, N711, N3182);
buf BUF1 (N4474, N4451);
and AND3 (N4475, N4467, N1286, N2938);
nor NOR4 (N4476, N4471, N3264, N1648, N4169);
nand NAND4 (N4477, N4475, N2139, N4360, N2138);
buf BUF1 (N4478, N4472);
buf BUF1 (N4479, N4465);
xor XOR2 (N4480, N4470, N4238);
xor XOR2 (N4481, N4477, N2645);
buf BUF1 (N4482, N4481);
not NOT1 (N4483, N4480);
nor NOR2 (N4484, N4482, N1039);
nor NOR3 (N4485, N4483, N3408, N969);
buf BUF1 (N4486, N4468);
not NOT1 (N4487, N4479);
nor NOR4 (N4488, N4487, N3075, N4325, N1069);
or OR2 (N4489, N4486, N638);
nor NOR3 (N4490, N4473, N4213, N1344);
xor XOR2 (N4491, N4474, N466);
buf BUF1 (N4492, N4478);
or OR4 (N4493, N4466, N2350, N1685, N4130);
nand NAND4 (N4494, N4489, N2308, N1036, N418);
buf BUF1 (N4495, N4488);
nor NOR3 (N4496, N4495, N3966, N3477);
nor NOR2 (N4497, N4490, N1954);
nor NOR2 (N4498, N4485, N3688);
nand NAND3 (N4499, N4436, N1605, N2334);
or OR2 (N4500, N4491, N3072);
xor XOR2 (N4501, N4497, N347);
nand NAND2 (N4502, N4484, N165);
and AND4 (N4503, N4502, N1771, N3693, N1381);
or OR2 (N4504, N4503, N3864);
not NOT1 (N4505, N4499);
buf BUF1 (N4506, N4505);
nor NOR2 (N4507, N4504, N1939);
nand NAND2 (N4508, N4494, N2428);
nor NOR3 (N4509, N4501, N292, N3734);
not NOT1 (N4510, N4500);
or OR2 (N4511, N4508, N1612);
nor NOR4 (N4512, N4509, N3029, N1006, N298);
nand NAND3 (N4513, N4506, N4300, N2846);
and AND3 (N4514, N4476, N2067, N1261);
not NOT1 (N4515, N4511);
and AND3 (N4516, N4498, N3041, N3627);
and AND3 (N4517, N4513, N2401, N3412);
and AND4 (N4518, N4514, N1938, N3044, N1621);
and AND4 (N4519, N4493, N3885, N777, N175);
nor NOR4 (N4520, N4517, N1437, N2281, N3792);
not NOT1 (N4521, N4519);
and AND4 (N4522, N4516, N2322, N3638, N3653);
not NOT1 (N4523, N4521);
not NOT1 (N4524, N4522);
or OR2 (N4525, N4496, N171);
not NOT1 (N4526, N4518);
and AND4 (N4527, N4515, N3127, N2653, N774);
nand NAND3 (N4528, N4520, N4183, N4047);
xor XOR2 (N4529, N4526, N4508);
buf BUF1 (N4530, N4507);
nand NAND4 (N4531, N4510, N2131, N2658, N2466);
nand NAND3 (N4532, N4529, N2517, N4405);
or OR4 (N4533, N4523, N2327, N3116, N1387);
xor XOR2 (N4534, N4512, N1397);
nor NOR4 (N4535, N4527, N759, N3933, N884);
or OR4 (N4536, N4533, N2232, N1881, N1193);
nand NAND2 (N4537, N4536, N1992);
nand NAND2 (N4538, N4524, N1515);
and AND3 (N4539, N4530, N4116, N2055);
not NOT1 (N4540, N4528);
xor XOR2 (N4541, N4534, N303);
or OR3 (N4542, N4532, N3418, N3183);
xor XOR2 (N4543, N4539, N417);
not NOT1 (N4544, N4492);
nand NAND4 (N4545, N4544, N1968, N1451, N1755);
nor NOR4 (N4546, N4542, N4467, N598, N3484);
or OR2 (N4547, N4531, N3129);
or OR3 (N4548, N4545, N735, N4405);
xor XOR2 (N4549, N4546, N2264);
xor XOR2 (N4550, N4538, N2965);
or OR2 (N4551, N4537, N2354);
nor NOR2 (N4552, N4540, N2529);
not NOT1 (N4553, N4543);
nand NAND2 (N4554, N4549, N1593);
buf BUF1 (N4555, N4535);
xor XOR2 (N4556, N4547, N2079);
not NOT1 (N4557, N4554);
and AND2 (N4558, N4557, N2977);
buf BUF1 (N4559, N4553);
or OR3 (N4560, N4541, N141, N492);
nand NAND2 (N4561, N4556, N529);
and AND2 (N4562, N4550, N1665);
buf BUF1 (N4563, N4558);
buf BUF1 (N4564, N4563);
buf BUF1 (N4565, N4552);
not NOT1 (N4566, N4561);
and AND3 (N4567, N4562, N2556, N2484);
xor XOR2 (N4568, N4567, N3910);
nor NOR4 (N4569, N4555, N2735, N4456, N4493);
nand NAND3 (N4570, N4560, N1873, N233);
buf BUF1 (N4571, N4551);
or OR3 (N4572, N4565, N4296, N1220);
and AND3 (N4573, N4559, N3334, N1153);
xor XOR2 (N4574, N4566, N3640);
nor NOR2 (N4575, N4564, N1905);
or OR4 (N4576, N4572, N3137, N106, N4553);
and AND2 (N4577, N4570, N82);
xor XOR2 (N4578, N4525, N925);
or OR4 (N4579, N4576, N4162, N1812, N2798);
buf BUF1 (N4580, N4578);
xor XOR2 (N4581, N4568, N909);
xor XOR2 (N4582, N4577, N3715);
nand NAND3 (N4583, N4571, N1367, N3314);
and AND3 (N4584, N4548, N278, N3817);
not NOT1 (N4585, N4569);
and AND3 (N4586, N4573, N4268, N2133);
or OR4 (N4587, N4580, N438, N1019, N2773);
nand NAND4 (N4588, N4587, N961, N85, N810);
and AND2 (N4589, N4574, N712);
xor XOR2 (N4590, N4586, N1947);
xor XOR2 (N4591, N4583, N1179);
nand NAND2 (N4592, N4584, N252);
nor NOR3 (N4593, N4581, N477, N1624);
xor XOR2 (N4594, N4588, N2178);
xor XOR2 (N4595, N4590, N3020);
or OR2 (N4596, N4594, N3064);
nor NOR2 (N4597, N4593, N184);
not NOT1 (N4598, N4589);
nand NAND2 (N4599, N4591, N4466);
and AND3 (N4600, N4592, N3948, N561);
and AND3 (N4601, N4596, N2269, N4215);
or OR4 (N4602, N4597, N2554, N605, N1430);
nand NAND2 (N4603, N4602, N4021);
xor XOR2 (N4604, N4582, N1178);
xor XOR2 (N4605, N4598, N206);
not NOT1 (N4606, N4575);
nor NOR2 (N4607, N4595, N3056);
not NOT1 (N4608, N4585);
or OR4 (N4609, N4579, N3369, N1360, N1598);
buf BUF1 (N4610, N4609);
nor NOR2 (N4611, N4608, N2040);
nand NAND3 (N4612, N4603, N3149, N1477);
nand NAND3 (N4613, N4599, N4347, N399);
nand NAND4 (N4614, N4600, N78, N1233, N2907);
or OR2 (N4615, N4606, N3620);
buf BUF1 (N4616, N4601);
buf BUF1 (N4617, N4611);
buf BUF1 (N4618, N4610);
nand NAND2 (N4619, N4605, N1605);
nor NOR2 (N4620, N4617, N2061);
and AND2 (N4621, N4620, N322);
nor NOR3 (N4622, N4615, N2405, N3280);
nand NAND3 (N4623, N4622, N4372, N2309);
and AND3 (N4624, N4618, N2718, N2672);
buf BUF1 (N4625, N4612);
nand NAND2 (N4626, N4614, N3488);
not NOT1 (N4627, N4613);
nor NOR4 (N4628, N4604, N679, N3452, N2166);
and AND2 (N4629, N4616, N3931);
xor XOR2 (N4630, N4626, N471);
buf BUF1 (N4631, N4628);
or OR4 (N4632, N4619, N1266, N4324, N1623);
buf BUF1 (N4633, N4632);
or OR4 (N4634, N4625, N2836, N1836, N3696);
nand NAND4 (N4635, N4623, N378, N808, N1626);
nor NOR2 (N4636, N4607, N3571);
or OR2 (N4637, N4634, N2177);
not NOT1 (N4638, N4631);
and AND3 (N4639, N4630, N374, N4338);
or OR4 (N4640, N4637, N3552, N1773, N2049);
xor XOR2 (N4641, N4638, N3552);
not NOT1 (N4642, N4639);
or OR4 (N4643, N4642, N4500, N2432, N4263);
nand NAND2 (N4644, N4643, N1426);
nor NOR3 (N4645, N4644, N1982, N4010);
nand NAND3 (N4646, N4629, N2738, N2537);
xor XOR2 (N4647, N4635, N4538);
or OR4 (N4648, N4647, N2185, N2818, N3963);
not NOT1 (N4649, N4627);
and AND4 (N4650, N4640, N3945, N56, N3170);
and AND2 (N4651, N4649, N275);
and AND4 (N4652, N4636, N650, N2124, N2977);
and AND2 (N4653, N4633, N2938);
buf BUF1 (N4654, N4651);
nor NOR4 (N4655, N4653, N2588, N326, N982);
nor NOR3 (N4656, N4650, N1328, N749);
nand NAND3 (N4657, N4621, N658, N2708);
xor XOR2 (N4658, N4655, N304);
or OR3 (N4659, N4654, N1232, N2214);
and AND2 (N4660, N4659, N2506);
xor XOR2 (N4661, N4646, N4127);
buf BUF1 (N4662, N4657);
not NOT1 (N4663, N4641);
or OR4 (N4664, N4656, N2318, N505, N4264);
and AND3 (N4665, N4664, N1852, N2845);
xor XOR2 (N4666, N4661, N4065);
buf BUF1 (N4667, N4645);
buf BUF1 (N4668, N4660);
buf BUF1 (N4669, N4668);
or OR4 (N4670, N4648, N3808, N2579, N2405);
xor XOR2 (N4671, N4663, N1568);
nand NAND2 (N4672, N4624, N1957);
xor XOR2 (N4673, N4666, N704);
xor XOR2 (N4674, N4671, N1014);
nor NOR3 (N4675, N4674, N4231, N4031);
and AND4 (N4676, N4665, N2488, N2208, N1916);
or OR4 (N4677, N4673, N3953, N3873, N4167);
or OR3 (N4678, N4675, N2410, N3668);
or OR2 (N4679, N4670, N2688);
and AND4 (N4680, N4677, N2528, N2497, N518);
and AND2 (N4681, N4667, N2174);
and AND3 (N4682, N4678, N4088, N615);
nor NOR2 (N4683, N4680, N3086);
not NOT1 (N4684, N4672);
and AND3 (N4685, N4683, N4555, N851);
not NOT1 (N4686, N4662);
nand NAND4 (N4687, N4682, N1749, N590, N4550);
xor XOR2 (N4688, N4679, N2478);
buf BUF1 (N4689, N4652);
nor NOR3 (N4690, N4686, N300, N2676);
or OR3 (N4691, N4676, N4069, N901);
buf BUF1 (N4692, N4691);
nor NOR3 (N4693, N4690, N3345, N392);
buf BUF1 (N4694, N4658);
or OR4 (N4695, N4692, N2432, N1743, N2933);
nor NOR3 (N4696, N4685, N1788, N2197);
or OR2 (N4697, N4684, N651);
buf BUF1 (N4698, N4669);
nor NOR4 (N4699, N4695, N3235, N2814, N417);
or OR2 (N4700, N4697, N4271);
not NOT1 (N4701, N4699);
not NOT1 (N4702, N4694);
and AND4 (N4703, N4687, N1266, N2109, N79);
or OR3 (N4704, N4696, N512, N1153);
not NOT1 (N4705, N4700);
or OR3 (N4706, N4688, N2943, N561);
or OR3 (N4707, N4706, N1510, N65);
nand NAND3 (N4708, N4701, N1485, N789);
and AND2 (N4709, N4705, N3084);
not NOT1 (N4710, N4704);
nor NOR2 (N4711, N4703, N3098);
buf BUF1 (N4712, N4708);
nor NOR2 (N4713, N4709, N2802);
and AND4 (N4714, N4689, N4119, N199, N3530);
or OR4 (N4715, N4681, N3999, N4045, N2090);
xor XOR2 (N4716, N4702, N2904);
nor NOR4 (N4717, N4715, N1664, N4085, N3165);
not NOT1 (N4718, N4711);
buf BUF1 (N4719, N4710);
xor XOR2 (N4720, N4712, N857);
not NOT1 (N4721, N4720);
xor XOR2 (N4722, N4693, N4458);
nor NOR2 (N4723, N4719, N3303);
nor NOR2 (N4724, N4717, N906);
buf BUF1 (N4725, N4718);
xor XOR2 (N4726, N4707, N1783);
buf BUF1 (N4727, N4723);
not NOT1 (N4728, N4726);
nor NOR4 (N4729, N4713, N4413, N1100, N829);
xor XOR2 (N4730, N4729, N2491);
or OR2 (N4731, N4721, N2118);
xor XOR2 (N4732, N4698, N2811);
or OR2 (N4733, N4727, N2180);
not NOT1 (N4734, N4722);
buf BUF1 (N4735, N4716);
buf BUF1 (N4736, N4725);
or OR2 (N4737, N4714, N3830);
nand NAND2 (N4738, N4724, N3999);
not NOT1 (N4739, N4737);
buf BUF1 (N4740, N4738);
nor NOR2 (N4741, N4739, N544);
or OR3 (N4742, N4740, N4071, N3019);
buf BUF1 (N4743, N4732);
or OR4 (N4744, N4730, N471, N86, N3458);
buf BUF1 (N4745, N4733);
buf BUF1 (N4746, N4743);
xor XOR2 (N4747, N4745, N3216);
or OR2 (N4748, N4731, N1992);
buf BUF1 (N4749, N4741);
nor NOR4 (N4750, N4749, N2223, N3962, N1558);
xor XOR2 (N4751, N4742, N162);
buf BUF1 (N4752, N4751);
nand NAND4 (N4753, N4750, N2586, N4123, N3107);
buf BUF1 (N4754, N4748);
buf BUF1 (N4755, N4747);
buf BUF1 (N4756, N4755);
and AND4 (N4757, N4746, N505, N2651, N3022);
nor NOR4 (N4758, N4756, N1541, N4241, N4338);
nand NAND2 (N4759, N4752, N219);
or OR3 (N4760, N4736, N946, N1407);
xor XOR2 (N4761, N4757, N819);
xor XOR2 (N4762, N4761, N3612);
buf BUF1 (N4763, N4762);
or OR2 (N4764, N4760, N2536);
nor NOR2 (N4765, N4764, N81);
buf BUF1 (N4766, N4765);
and AND3 (N4767, N4728, N1604, N1828);
or OR2 (N4768, N4734, N555);
not NOT1 (N4769, N4767);
nor NOR2 (N4770, N4769, N1906);
nand NAND3 (N4771, N4770, N3735, N3797);
and AND4 (N4772, N4744, N1732, N3353, N2887);
or OR3 (N4773, N4754, N3741, N1829);
or OR3 (N4774, N4758, N766, N616);
xor XOR2 (N4775, N4771, N3352);
xor XOR2 (N4776, N4753, N687);
or OR2 (N4777, N4776, N1376);
not NOT1 (N4778, N4773);
buf BUF1 (N4779, N4735);
not NOT1 (N4780, N4772);
or OR3 (N4781, N4774, N4361, N217);
and AND4 (N4782, N4779, N3604, N3366, N2972);
or OR3 (N4783, N4777, N2442, N862);
or OR3 (N4784, N4780, N4118, N2242);
xor XOR2 (N4785, N4784, N2683);
not NOT1 (N4786, N4778);
nand NAND3 (N4787, N4766, N403, N1052);
buf BUF1 (N4788, N4781);
nor NOR4 (N4789, N4775, N3461, N4619, N3483);
and AND3 (N4790, N4783, N373, N1756);
nand NAND3 (N4791, N4763, N2906, N1283);
not NOT1 (N4792, N4786);
and AND3 (N4793, N4789, N838, N2978);
nor NOR3 (N4794, N4788, N3762, N4234);
nor NOR3 (N4795, N4791, N1161, N4276);
not NOT1 (N4796, N4795);
nand NAND3 (N4797, N4790, N519, N2691);
and AND2 (N4798, N4794, N105);
or OR2 (N4799, N4793, N1380);
buf BUF1 (N4800, N4798);
and AND2 (N4801, N4796, N1249);
buf BUF1 (N4802, N4801);
buf BUF1 (N4803, N4782);
xor XOR2 (N4804, N4800, N1643);
and AND4 (N4805, N4759, N2248, N4560, N3613);
buf BUF1 (N4806, N4799);
nor NOR2 (N4807, N4797, N2800);
nand NAND3 (N4808, N4807, N2889, N4775);
buf BUF1 (N4809, N4806);
or OR2 (N4810, N4804, N4792);
not NOT1 (N4811, N98);
or OR3 (N4812, N4809, N4431, N3498);
buf BUF1 (N4813, N4787);
or OR2 (N4814, N4802, N2463);
not NOT1 (N4815, N4810);
nor NOR2 (N4816, N4814, N1815);
xor XOR2 (N4817, N4808, N1149);
buf BUF1 (N4818, N4805);
not NOT1 (N4819, N4816);
not NOT1 (N4820, N4817);
not NOT1 (N4821, N4812);
xor XOR2 (N4822, N4821, N2220);
or OR2 (N4823, N4820, N1924);
nor NOR3 (N4824, N4818, N2149, N370);
nor NOR2 (N4825, N4824, N2807);
and AND2 (N4826, N4803, N443);
nand NAND4 (N4827, N4826, N2131, N2482, N4092);
nand NAND3 (N4828, N4815, N3635, N3621);
nand NAND2 (N4829, N4828, N2114);
or OR4 (N4830, N4823, N4068, N3100, N4474);
or OR3 (N4831, N4811, N3724, N1972);
or OR2 (N4832, N4813, N1455);
nand NAND3 (N4833, N4831, N2097, N97);
and AND3 (N4834, N4785, N1817, N77);
xor XOR2 (N4835, N4825, N1749);
or OR3 (N4836, N4832, N321, N3866);
nor NOR3 (N4837, N4827, N20, N4266);
not NOT1 (N4838, N4768);
nand NAND3 (N4839, N4829, N2461, N4508);
not NOT1 (N4840, N4819);
and AND4 (N4841, N4839, N4099, N3166, N3364);
xor XOR2 (N4842, N4841, N3658);
buf BUF1 (N4843, N4833);
xor XOR2 (N4844, N4837, N3168);
not NOT1 (N4845, N4844);
or OR2 (N4846, N4834, N286);
and AND4 (N4847, N4835, N421, N636, N297);
not NOT1 (N4848, N4822);
or OR2 (N4849, N4836, N3635);
buf BUF1 (N4850, N4847);
and AND4 (N4851, N4840, N2468, N2864, N2474);
nor NOR3 (N4852, N4838, N2451, N1070);
nand NAND3 (N4853, N4845, N4368, N3574);
not NOT1 (N4854, N4852);
and AND2 (N4855, N4848, N2711);
not NOT1 (N4856, N4849);
nor NOR2 (N4857, N4830, N4758);
not NOT1 (N4858, N4842);
nor NOR4 (N4859, N4843, N3503, N4568, N2035);
and AND3 (N4860, N4857, N64, N693);
or OR2 (N4861, N4850, N2494);
xor XOR2 (N4862, N4860, N1893);
nor NOR2 (N4863, N4853, N750);
nor NOR2 (N4864, N4861, N595);
buf BUF1 (N4865, N4863);
or OR4 (N4866, N4854, N3899, N1642, N3710);
buf BUF1 (N4867, N4859);
buf BUF1 (N4868, N4856);
or OR4 (N4869, N4866, N823, N659, N429);
nand NAND4 (N4870, N4855, N4763, N682, N4488);
xor XOR2 (N4871, N4858, N835);
or OR3 (N4872, N4865, N1189, N3542);
nand NAND3 (N4873, N4867, N3809, N2222);
and AND3 (N4874, N4868, N3003, N3076);
xor XOR2 (N4875, N4870, N3898);
not NOT1 (N4876, N4869);
or OR2 (N4877, N4846, N2994);
buf BUF1 (N4878, N4862);
nor NOR4 (N4879, N4877, N573, N3297, N4208);
buf BUF1 (N4880, N4878);
xor XOR2 (N4881, N4851, N2267);
and AND2 (N4882, N4881, N3964);
nor NOR3 (N4883, N4874, N3914, N719);
and AND4 (N4884, N4879, N4168, N2341, N1862);
nor NOR3 (N4885, N4884, N1812, N337);
nand NAND3 (N4886, N4873, N3292, N3649);
nand NAND4 (N4887, N4885, N2538, N2163, N3257);
nand NAND4 (N4888, N4880, N2954, N1035, N2239);
nor NOR3 (N4889, N4888, N2493, N1754);
buf BUF1 (N4890, N4887);
and AND2 (N4891, N4864, N3224);
xor XOR2 (N4892, N4882, N4286);
nor NOR2 (N4893, N4890, N4757);
and AND2 (N4894, N4871, N575);
and AND4 (N4895, N4883, N3104, N4558, N1946);
nor NOR4 (N4896, N4891, N2682, N3112, N2820);
and AND3 (N4897, N4893, N3759, N3307);
or OR2 (N4898, N4892, N302);
not NOT1 (N4899, N4875);
xor XOR2 (N4900, N4896, N1104);
xor XOR2 (N4901, N4886, N438);
or OR4 (N4902, N4901, N4051, N3185, N3698);
nor NOR2 (N4903, N4889, N1471);
or OR4 (N4904, N4895, N2626, N3332, N975);
or OR4 (N4905, N4903, N3965, N2082, N3051);
and AND3 (N4906, N4894, N2450, N2215);
not NOT1 (N4907, N4898);
buf BUF1 (N4908, N4900);
not NOT1 (N4909, N4897);
not NOT1 (N4910, N4904);
nand NAND4 (N4911, N4876, N853, N1089, N3040);
nand NAND4 (N4912, N4911, N4183, N3400, N4271);
or OR4 (N4913, N4905, N4495, N2310, N951);
nand NAND3 (N4914, N4902, N2741, N300);
nand NAND4 (N4915, N4907, N895, N4486, N990);
or OR3 (N4916, N4908, N3531, N3105);
not NOT1 (N4917, N4914);
nor NOR2 (N4918, N4910, N3721);
buf BUF1 (N4919, N4909);
nor NOR2 (N4920, N4918, N1120);
xor XOR2 (N4921, N4913, N3552);
and AND2 (N4922, N4916, N3372);
or OR3 (N4923, N4917, N1764, N801);
not NOT1 (N4924, N4921);
and AND3 (N4925, N4915, N379, N4274);
xor XOR2 (N4926, N4906, N984);
nor NOR2 (N4927, N4920, N180);
buf BUF1 (N4928, N4922);
nand NAND2 (N4929, N4923, N2567);
buf BUF1 (N4930, N4927);
and AND2 (N4931, N4929, N1288);
nor NOR3 (N4932, N4872, N1355, N4457);
xor XOR2 (N4933, N4926, N674);
nor NOR2 (N4934, N4928, N1929);
or OR4 (N4935, N4899, N371, N4233, N504);
buf BUF1 (N4936, N4930);
xor XOR2 (N4937, N4919, N3954);
buf BUF1 (N4938, N4925);
nand NAND4 (N4939, N4936, N989, N3557, N1214);
xor XOR2 (N4940, N4938, N100);
xor XOR2 (N4941, N4934, N120);
nand NAND2 (N4942, N4932, N3924);
xor XOR2 (N4943, N4924, N3383);
buf BUF1 (N4944, N4933);
and AND2 (N4945, N4944, N383);
not NOT1 (N4946, N4941);
nor NOR2 (N4947, N4937, N501);
nor NOR2 (N4948, N4939, N4367);
and AND2 (N4949, N4940, N697);
nor NOR3 (N4950, N4945, N2467, N2482);
xor XOR2 (N4951, N4950, N1774);
xor XOR2 (N4952, N4942, N157);
and AND3 (N4953, N4912, N1672, N1356);
and AND2 (N4954, N4949, N570);
nand NAND4 (N4955, N4951, N2057, N3417, N2865);
or OR2 (N4956, N4952, N407);
xor XOR2 (N4957, N4947, N1420);
buf BUF1 (N4958, N4953);
not NOT1 (N4959, N4943);
nor NOR3 (N4960, N4958, N1952, N2546);
not NOT1 (N4961, N4956);
xor XOR2 (N4962, N4960, N2644);
or OR2 (N4963, N4948, N1188);
nand NAND4 (N4964, N4955, N1107, N334, N4907);
xor XOR2 (N4965, N4961, N4935);
nand NAND2 (N4966, N513, N2614);
not NOT1 (N4967, N4959);
nand NAND4 (N4968, N4954, N3014, N3012, N2844);
and AND4 (N4969, N4946, N3314, N1652, N737);
or OR2 (N4970, N4968, N3603);
xor XOR2 (N4971, N4967, N905);
nand NAND3 (N4972, N4971, N2851, N3528);
not NOT1 (N4973, N4931);
xor XOR2 (N4974, N4969, N870);
nor NOR2 (N4975, N4957, N1038);
or OR3 (N4976, N4963, N1809, N877);
not NOT1 (N4977, N4962);
buf BUF1 (N4978, N4977);
and AND4 (N4979, N4970, N1782, N1576, N3954);
nor NOR4 (N4980, N4972, N2442, N4474, N4086);
xor XOR2 (N4981, N4974, N2947);
and AND2 (N4982, N4978, N4256);
and AND2 (N4983, N4981, N4388);
not NOT1 (N4984, N4983);
not NOT1 (N4985, N4976);
nand NAND3 (N4986, N4964, N1909, N1957);
nand NAND2 (N4987, N4985, N2791);
nand NAND3 (N4988, N4965, N1687, N4919);
not NOT1 (N4989, N4979);
buf BUF1 (N4990, N4987);
not NOT1 (N4991, N4989);
xor XOR2 (N4992, N4975, N4415);
not NOT1 (N4993, N4973);
nor NOR2 (N4994, N4986, N3949);
and AND4 (N4995, N4988, N3339, N4007, N1162);
and AND3 (N4996, N4980, N475, N3739);
xor XOR2 (N4997, N4991, N328);
and AND3 (N4998, N4982, N1120, N1396);
nor NOR2 (N4999, N4984, N3694);
and AND4 (N5000, N4994, N1910, N4417, N4189);
or OR3 (N5001, N4996, N4354, N1630);
and AND3 (N5002, N4997, N79, N4053);
nor NOR4 (N5003, N4966, N4359, N2243, N975);
xor XOR2 (N5004, N4990, N3395);
nor NOR3 (N5005, N4992, N4853, N1856);
xor XOR2 (N5006, N5003, N1412);
nand NAND4 (N5007, N4999, N629, N3100, N4275);
nand NAND2 (N5008, N4998, N3959);
xor XOR2 (N5009, N5005, N848);
and AND2 (N5010, N5006, N4667);
nor NOR4 (N5011, N4993, N4006, N3690, N17);
buf BUF1 (N5012, N5009);
and AND4 (N5013, N5010, N534, N415, N52);
not NOT1 (N5014, N5004);
buf BUF1 (N5015, N5001);
not NOT1 (N5016, N5015);
buf BUF1 (N5017, N5002);
xor XOR2 (N5018, N5016, N598);
not NOT1 (N5019, N5012);
xor XOR2 (N5020, N5018, N2989);
or OR3 (N5021, N5013, N4502, N2043);
not NOT1 (N5022, N5011);
and AND3 (N5023, N5021, N1496, N438);
or OR3 (N5024, N5007, N4116, N513);
or OR2 (N5025, N5014, N2467);
nor NOR4 (N5026, N5017, N1398, N4734, N1559);
buf BUF1 (N5027, N5008);
and AND2 (N5028, N4995, N3922);
and AND4 (N5029, N5026, N226, N1995, N2737);
nand NAND4 (N5030, N5029, N3170, N323, N4363);
or OR4 (N5031, N5028, N1676, N4235, N5005);
buf BUF1 (N5032, N5019);
and AND2 (N5033, N5023, N3622);
nand NAND2 (N5034, N5000, N433);
and AND2 (N5035, N5034, N2871);
or OR2 (N5036, N5025, N3265);
and AND3 (N5037, N5020, N2815, N1920);
xor XOR2 (N5038, N5032, N683);
or OR4 (N5039, N5024, N464, N4829, N3567);
not NOT1 (N5040, N5033);
or OR2 (N5041, N5037, N3499);
buf BUF1 (N5042, N5031);
nor NOR3 (N5043, N5027, N1921, N247);
nand NAND2 (N5044, N5043, N94);
xor XOR2 (N5045, N5044, N1120);
nand NAND3 (N5046, N5022, N4863, N914);
buf BUF1 (N5047, N5041);
and AND3 (N5048, N5040, N2719, N2484);
or OR2 (N5049, N5035, N628);
xor XOR2 (N5050, N5038, N4818);
buf BUF1 (N5051, N5030);
not NOT1 (N5052, N5039);
or OR2 (N5053, N5042, N3806);
and AND2 (N5054, N5052, N4996);
not NOT1 (N5055, N5046);
and AND2 (N5056, N5048, N683);
or OR4 (N5057, N5056, N2810, N221, N46);
nor NOR2 (N5058, N5057, N1489);
or OR3 (N5059, N5058, N1087, N1730);
xor XOR2 (N5060, N5049, N4425);
not NOT1 (N5061, N5059);
not NOT1 (N5062, N5036);
buf BUF1 (N5063, N5045);
and AND4 (N5064, N5051, N354, N706, N384);
and AND4 (N5065, N5054, N2116, N4056, N2527);
nor NOR4 (N5066, N5064, N3885, N4002, N3846);
xor XOR2 (N5067, N5050, N3170);
not NOT1 (N5068, N5055);
xor XOR2 (N5069, N5063, N276);
buf BUF1 (N5070, N5065);
or OR3 (N5071, N5062, N4926, N3079);
or OR4 (N5072, N5047, N3106, N2656, N203);
nor NOR3 (N5073, N5069, N494, N1779);
xor XOR2 (N5074, N5061, N451);
or OR2 (N5075, N5068, N3902);
not NOT1 (N5076, N5074);
and AND3 (N5077, N5075, N925, N3658);
xor XOR2 (N5078, N5067, N5003);
buf BUF1 (N5079, N5060);
buf BUF1 (N5080, N5078);
nor NOR4 (N5081, N5071, N1959, N2501, N1);
or OR3 (N5082, N5073, N2333, N2277);
not NOT1 (N5083, N5079);
nand NAND4 (N5084, N5083, N2841, N4787, N999);
or OR4 (N5085, N5082, N1940, N4026, N4280);
and AND4 (N5086, N5085, N840, N1095, N4114);
xor XOR2 (N5087, N5077, N4228);
nand NAND4 (N5088, N5072, N2068, N2061, N3565);
and AND3 (N5089, N5088, N681, N2190);
xor XOR2 (N5090, N5070, N1740);
and AND2 (N5091, N5090, N1445);
nand NAND3 (N5092, N5053, N3225, N3709);
or OR2 (N5093, N5081, N2565);
or OR2 (N5094, N5086, N1893);
not NOT1 (N5095, N5087);
nand NAND2 (N5096, N5089, N1922);
and AND3 (N5097, N5093, N1991, N298);
not NOT1 (N5098, N5095);
and AND2 (N5099, N5076, N188);
or OR4 (N5100, N5066, N3156, N2674, N3724);
or OR4 (N5101, N5080, N1344, N3354, N1134);
nand NAND4 (N5102, N5098, N444, N3877, N845);
and AND2 (N5103, N5096, N2955);
buf BUF1 (N5104, N5103);
nand NAND2 (N5105, N5091, N138);
not NOT1 (N5106, N5101);
nor NOR2 (N5107, N5092, N2709);
nand NAND2 (N5108, N5084, N746);
or OR2 (N5109, N5106, N858);
not NOT1 (N5110, N5094);
or OR3 (N5111, N5110, N4112, N1714);
and AND2 (N5112, N5099, N526);
not NOT1 (N5113, N5104);
buf BUF1 (N5114, N5111);
or OR2 (N5115, N5108, N3234);
nand NAND2 (N5116, N5113, N779);
xor XOR2 (N5117, N5107, N2002);
nor NOR4 (N5118, N5109, N3232, N1223, N4929);
xor XOR2 (N5119, N5115, N188);
or OR3 (N5120, N5112, N806, N2691);
not NOT1 (N5121, N5102);
xor XOR2 (N5122, N5120, N2710);
nor NOR3 (N5123, N5122, N3142, N4510);
nor NOR2 (N5124, N5116, N4656);
nor NOR3 (N5125, N5119, N4379, N144);
or OR4 (N5126, N5118, N2791, N2388, N517);
and AND4 (N5127, N5105, N4631, N2269, N4717);
or OR3 (N5128, N5097, N2116, N2781);
nor NOR4 (N5129, N5125, N3649, N2275, N109);
buf BUF1 (N5130, N5124);
not NOT1 (N5131, N5114);
xor XOR2 (N5132, N5126, N4501);
not NOT1 (N5133, N5127);
not NOT1 (N5134, N5121);
buf BUF1 (N5135, N5133);
and AND4 (N5136, N5130, N1279, N555, N3411);
or OR3 (N5137, N5129, N2677, N2952);
and AND4 (N5138, N5131, N1804, N5123, N2928);
xor XOR2 (N5139, N4888, N2851);
not NOT1 (N5140, N5135);
or OR4 (N5141, N5140, N3586, N510, N687);
not NOT1 (N5142, N5141);
or OR3 (N5143, N5138, N3328, N1161);
nand NAND3 (N5144, N5117, N3809, N1448);
or OR2 (N5145, N5134, N110);
nor NOR4 (N5146, N5100, N1359, N3116, N3142);
xor XOR2 (N5147, N5142, N1826);
xor XOR2 (N5148, N5143, N4709);
or OR4 (N5149, N5136, N4728, N4619, N2922);
or OR4 (N5150, N5147, N905, N3633, N814);
nand NAND3 (N5151, N5137, N3861, N2656);
xor XOR2 (N5152, N5145, N1290);
nor NOR4 (N5153, N5151, N376, N1648, N1473);
and AND4 (N5154, N5139, N727, N675, N1174);
xor XOR2 (N5155, N5128, N1930);
not NOT1 (N5156, N5150);
nor NOR3 (N5157, N5156, N2096, N1533);
nand NAND2 (N5158, N5157, N740);
nor NOR3 (N5159, N5154, N5115, N2140);
not NOT1 (N5160, N5152);
not NOT1 (N5161, N5148);
nor NOR4 (N5162, N5161, N1833, N5100, N318);
nand NAND3 (N5163, N5149, N433, N2273);
not NOT1 (N5164, N5160);
and AND2 (N5165, N5164, N1047);
nor NOR2 (N5166, N5155, N1174);
nand NAND2 (N5167, N5163, N405);
and AND3 (N5168, N5158, N807, N2596);
nor NOR3 (N5169, N5159, N979, N388);
xor XOR2 (N5170, N5166, N2852);
xor XOR2 (N5171, N5165, N1575);
xor XOR2 (N5172, N5153, N2041);
and AND2 (N5173, N5172, N3719);
or OR2 (N5174, N5167, N188);
or OR4 (N5175, N5169, N4369, N3199, N2497);
nand NAND2 (N5176, N5162, N5155);
and AND2 (N5177, N5144, N4448);
not NOT1 (N5178, N5170);
buf BUF1 (N5179, N5146);
or OR2 (N5180, N5175, N1242);
nand NAND4 (N5181, N5178, N2749, N1528, N2096);
not NOT1 (N5182, N5171);
nand NAND3 (N5183, N5173, N3167, N4004);
or OR3 (N5184, N5177, N5162, N5057);
nor NOR2 (N5185, N5183, N3636);
nor NOR2 (N5186, N5182, N2570);
nor NOR4 (N5187, N5184, N1327, N4401, N4140);
nand NAND3 (N5188, N5176, N2357, N1066);
or OR2 (N5189, N5188, N2593);
nand NAND3 (N5190, N5174, N3360, N3789);
nand NAND2 (N5191, N5185, N3475);
nor NOR3 (N5192, N5187, N4943, N2537);
xor XOR2 (N5193, N5179, N1653);
nor NOR2 (N5194, N5180, N32);
buf BUF1 (N5195, N5192);
nand NAND2 (N5196, N5168, N1882);
or OR2 (N5197, N5190, N4599);
not NOT1 (N5198, N5181);
nand NAND2 (N5199, N5132, N4774);
or OR2 (N5200, N5193, N1164);
nor NOR2 (N5201, N5196, N832);
nand NAND2 (N5202, N5199, N2620);
or OR2 (N5203, N5200, N510);
nand NAND3 (N5204, N5201, N2747, N4987);
and AND3 (N5205, N5194, N2265, N3593);
and AND3 (N5206, N5195, N4224, N2589);
not NOT1 (N5207, N5205);
buf BUF1 (N5208, N5191);
not NOT1 (N5209, N5207);
and AND4 (N5210, N5189, N4593, N3458, N608);
buf BUF1 (N5211, N5186);
and AND2 (N5212, N5202, N2053);
buf BUF1 (N5213, N5209);
or OR2 (N5214, N5210, N2964);
buf BUF1 (N5215, N5211);
and AND3 (N5216, N5198, N484, N4616);
and AND4 (N5217, N5197, N1673, N213, N3436);
nor NOR4 (N5218, N5217, N1221, N2936, N1144);
xor XOR2 (N5219, N5213, N3820);
nor NOR3 (N5220, N5216, N5137, N4427);
not NOT1 (N5221, N5208);
buf BUF1 (N5222, N5220);
not NOT1 (N5223, N5206);
nand NAND4 (N5224, N5223, N2612, N1816, N321);
not NOT1 (N5225, N5215);
and AND4 (N5226, N5212, N1519, N2038, N1330);
buf BUF1 (N5227, N5204);
or OR4 (N5228, N5226, N3812, N1655, N187);
not NOT1 (N5229, N5214);
and AND2 (N5230, N5222, N1193);
and AND2 (N5231, N5224, N2651);
and AND4 (N5232, N5218, N4123, N1218, N493);
xor XOR2 (N5233, N5221, N4013);
buf BUF1 (N5234, N5225);
and AND3 (N5235, N5228, N1432, N5010);
nand NAND3 (N5236, N5231, N5148, N1183);
nor NOR4 (N5237, N5219, N2614, N2402, N3625);
or OR2 (N5238, N5230, N139);
or OR2 (N5239, N5235, N435);
nor NOR3 (N5240, N5203, N1710, N296);
or OR4 (N5241, N5236, N4971, N369, N1793);
not NOT1 (N5242, N5238);
xor XOR2 (N5243, N5237, N2729);
or OR2 (N5244, N5239, N2218);
xor XOR2 (N5245, N5227, N4143);
xor XOR2 (N5246, N5229, N1593);
or OR4 (N5247, N5241, N4449, N2385, N3257);
nand NAND4 (N5248, N5246, N508, N3880, N4504);
and AND4 (N5249, N5248, N1933, N2131, N2230);
xor XOR2 (N5250, N5245, N3702);
or OR3 (N5251, N5234, N5214, N5099);
and AND4 (N5252, N5249, N4170, N497, N4008);
nor NOR3 (N5253, N5243, N3223, N1739);
xor XOR2 (N5254, N5251, N614);
or OR3 (N5255, N5252, N4572, N3998);
xor XOR2 (N5256, N5253, N5247);
or OR2 (N5257, N5239, N3925);
and AND2 (N5258, N5244, N2787);
nand NAND4 (N5259, N5240, N998, N4284, N334);
nor NOR3 (N5260, N5242, N3973, N4857);
xor XOR2 (N5261, N5250, N1358);
buf BUF1 (N5262, N5257);
and AND2 (N5263, N5261, N4089);
not NOT1 (N5264, N5263);
or OR3 (N5265, N5256, N854, N2174);
xor XOR2 (N5266, N5264, N4969);
xor XOR2 (N5267, N5265, N65);
and AND4 (N5268, N5254, N2232, N100, N751);
buf BUF1 (N5269, N5266);
and AND4 (N5270, N5258, N5134, N3097, N986);
or OR4 (N5271, N5262, N4095, N1521, N3407);
buf BUF1 (N5272, N5267);
not NOT1 (N5273, N5259);
or OR4 (N5274, N5232, N2006, N5125, N4271);
nor NOR2 (N5275, N5270, N2552);
buf BUF1 (N5276, N5268);
and AND4 (N5277, N5272, N1437, N5275, N37);
not NOT1 (N5278, N3292);
not NOT1 (N5279, N5255);
and AND3 (N5280, N5269, N683, N2844);
buf BUF1 (N5281, N5273);
xor XOR2 (N5282, N5276, N1228);
not NOT1 (N5283, N5280);
and AND2 (N5284, N5279, N2912);
and AND4 (N5285, N5284, N875, N1501, N2802);
nor NOR3 (N5286, N5274, N841, N4463);
not NOT1 (N5287, N5278);
nand NAND4 (N5288, N5283, N2265, N1670, N4725);
and AND2 (N5289, N5286, N1018);
and AND2 (N5290, N5233, N36);
xor XOR2 (N5291, N5288, N1954);
buf BUF1 (N5292, N5289);
xor XOR2 (N5293, N5287, N5277);
buf BUF1 (N5294, N574);
not NOT1 (N5295, N5285);
nand NAND4 (N5296, N5292, N5182, N5231, N14);
nor NOR2 (N5297, N5290, N2273);
nor NOR2 (N5298, N5294, N2690);
buf BUF1 (N5299, N5291);
and AND2 (N5300, N5297, N911);
and AND2 (N5301, N5300, N922);
xor XOR2 (N5302, N5295, N3613);
nor NOR3 (N5303, N5299, N869, N1869);
not NOT1 (N5304, N5293);
and AND2 (N5305, N5296, N3561);
xor XOR2 (N5306, N5281, N1729);
xor XOR2 (N5307, N5298, N4390);
or OR3 (N5308, N5282, N1769, N4507);
buf BUF1 (N5309, N5301);
and AND4 (N5310, N5305, N1843, N666, N3435);
nand NAND2 (N5311, N5304, N494);
not NOT1 (N5312, N5311);
not NOT1 (N5313, N5260);
xor XOR2 (N5314, N5302, N1124);
and AND4 (N5315, N5271, N1927, N4484, N3472);
nand NAND2 (N5316, N5314, N2641);
nand NAND2 (N5317, N5310, N665);
and AND4 (N5318, N5309, N4722, N2137, N1138);
xor XOR2 (N5319, N5303, N2655);
nand NAND4 (N5320, N5315, N2266, N1091, N3154);
nor NOR4 (N5321, N5307, N1593, N2515, N3272);
not NOT1 (N5322, N5317);
nor NOR3 (N5323, N5320, N4316, N2607);
and AND3 (N5324, N5321, N2090, N4562);
xor XOR2 (N5325, N5308, N3191);
nor NOR4 (N5326, N5306, N4675, N1097, N2000);
nand NAND4 (N5327, N5319, N3501, N65, N2631);
buf BUF1 (N5328, N5326);
buf BUF1 (N5329, N5312);
nand NAND2 (N5330, N5323, N2810);
nor NOR3 (N5331, N5325, N295, N4317);
xor XOR2 (N5332, N5318, N4909);
buf BUF1 (N5333, N5322);
not NOT1 (N5334, N5331);
not NOT1 (N5335, N5316);
nand NAND2 (N5336, N5328, N4791);
not NOT1 (N5337, N5329);
xor XOR2 (N5338, N5333, N1835);
buf BUF1 (N5339, N5313);
or OR4 (N5340, N5332, N5206, N5080, N4196);
or OR2 (N5341, N5335, N2509);
and AND3 (N5342, N5338, N2759, N291);
xor XOR2 (N5343, N5342, N747);
nor NOR3 (N5344, N5327, N3511, N503);
not NOT1 (N5345, N5340);
nor NOR3 (N5346, N5344, N2125, N963);
nand NAND3 (N5347, N5341, N1951, N3218);
buf BUF1 (N5348, N5343);
xor XOR2 (N5349, N5346, N2595);
nand NAND4 (N5350, N5348, N4162, N2185, N3870);
or OR3 (N5351, N5334, N2944, N3359);
buf BUF1 (N5352, N5349);
and AND2 (N5353, N5324, N3563);
nor NOR3 (N5354, N5336, N4298, N1281);
or OR3 (N5355, N5337, N4049, N5256);
buf BUF1 (N5356, N5330);
buf BUF1 (N5357, N5355);
xor XOR2 (N5358, N5345, N1818);
or OR4 (N5359, N5356, N4397, N1302, N1393);
and AND3 (N5360, N5350, N1691, N1823);
nor NOR4 (N5361, N5347, N1829, N93, N4432);
and AND2 (N5362, N5360, N4451);
buf BUF1 (N5363, N5359);
or OR2 (N5364, N5362, N57);
not NOT1 (N5365, N5354);
nor NOR4 (N5366, N5361, N2072, N43, N5205);
nand NAND2 (N5367, N5351, N3760);
not NOT1 (N5368, N5357);
nor NOR2 (N5369, N5358, N2117);
xor XOR2 (N5370, N5364, N2449);
buf BUF1 (N5371, N5352);
buf BUF1 (N5372, N5366);
nand NAND3 (N5373, N5369, N2430, N3318);
xor XOR2 (N5374, N5365, N4620);
not NOT1 (N5375, N5339);
xor XOR2 (N5376, N5371, N2607);
xor XOR2 (N5377, N5363, N84);
xor XOR2 (N5378, N5374, N2860);
xor XOR2 (N5379, N5370, N1980);
buf BUF1 (N5380, N5372);
and AND4 (N5381, N5379, N5158, N3054, N3417);
nor NOR3 (N5382, N5380, N2107, N4692);
or OR3 (N5383, N5368, N4113, N1237);
nor NOR4 (N5384, N5378, N4195, N1553, N2946);
not NOT1 (N5385, N5384);
or OR4 (N5386, N5377, N4506, N4679, N815);
not NOT1 (N5387, N5375);
nand NAND3 (N5388, N5386, N1073, N4365);
nand NAND2 (N5389, N5382, N366);
not NOT1 (N5390, N5383);
or OR4 (N5391, N5390, N3797, N5331, N1097);
xor XOR2 (N5392, N5388, N940);
buf BUF1 (N5393, N5387);
nand NAND4 (N5394, N5376, N3092, N370, N4657);
and AND2 (N5395, N5367, N4297);
not NOT1 (N5396, N5353);
buf BUF1 (N5397, N5394);
buf BUF1 (N5398, N5389);
and AND2 (N5399, N5396, N4767);
and AND4 (N5400, N5381, N970, N1313, N4933);
nand NAND2 (N5401, N5397, N2607);
or OR3 (N5402, N5393, N5206, N4908);
xor XOR2 (N5403, N5398, N723);
or OR2 (N5404, N5400, N5189);
nand NAND3 (N5405, N5385, N1349, N1510);
and AND3 (N5406, N5395, N3790, N3496);
buf BUF1 (N5407, N5403);
xor XOR2 (N5408, N5402, N3963);
xor XOR2 (N5409, N5391, N1676);
nand NAND2 (N5410, N5401, N4810);
or OR3 (N5411, N5392, N4602, N492);
nor NOR3 (N5412, N5373, N1886, N4426);
not NOT1 (N5413, N5411);
nor NOR4 (N5414, N5407, N1792, N4505, N4685);
nand NAND3 (N5415, N5409, N3904, N4352);
and AND3 (N5416, N5404, N1098, N2824);
nor NOR2 (N5417, N5399, N532);
buf BUF1 (N5418, N5414);
buf BUF1 (N5419, N5412);
buf BUF1 (N5420, N5405);
buf BUF1 (N5421, N5408);
xor XOR2 (N5422, N5420, N192);
or OR4 (N5423, N5417, N2419, N3041, N3444);
nand NAND2 (N5424, N5410, N5079);
xor XOR2 (N5425, N5421, N4687);
or OR2 (N5426, N5424, N5103);
xor XOR2 (N5427, N5413, N1259);
not NOT1 (N5428, N5419);
or OR3 (N5429, N5416, N1046, N552);
not NOT1 (N5430, N5428);
or OR2 (N5431, N5415, N4758);
nor NOR2 (N5432, N5418, N423);
nor NOR2 (N5433, N5429, N296);
and AND2 (N5434, N5431, N5005);
not NOT1 (N5435, N5434);
and AND3 (N5436, N5435, N1066, N504);
nand NAND2 (N5437, N5427, N638);
nand NAND3 (N5438, N5433, N3171, N3300);
nor NOR3 (N5439, N5422, N2611, N2759);
buf BUF1 (N5440, N5437);
nand NAND3 (N5441, N5438, N3501, N650);
xor XOR2 (N5442, N5406, N1770);
xor XOR2 (N5443, N5425, N4091);
buf BUF1 (N5444, N5441);
or OR3 (N5445, N5423, N4234, N3360);
xor XOR2 (N5446, N5430, N4510);
buf BUF1 (N5447, N5443);
xor XOR2 (N5448, N5444, N5399);
or OR2 (N5449, N5432, N297);
not NOT1 (N5450, N5446);
xor XOR2 (N5451, N5449, N281);
or OR4 (N5452, N5448, N862, N5061, N661);
nor NOR2 (N5453, N5450, N3016);
not NOT1 (N5454, N5453);
nand NAND4 (N5455, N5440, N1931, N2906, N615);
not NOT1 (N5456, N5439);
nand NAND2 (N5457, N5442, N1053);
nand NAND2 (N5458, N5447, N3713);
buf BUF1 (N5459, N5455);
nand NAND4 (N5460, N5451, N1720, N3144, N690);
nand NAND2 (N5461, N5452, N4485);
not NOT1 (N5462, N5426);
and AND2 (N5463, N5460, N186);
xor XOR2 (N5464, N5461, N4704);
nand NAND4 (N5465, N5436, N4502, N2489, N2413);
and AND2 (N5466, N5445, N3819);
buf BUF1 (N5467, N5465);
xor XOR2 (N5468, N5457, N672);
nor NOR2 (N5469, N5458, N3518);
and AND4 (N5470, N5459, N492, N1881, N4121);
xor XOR2 (N5471, N5464, N1613);
nand NAND2 (N5472, N5456, N5371);
nand NAND4 (N5473, N5468, N2127, N2173, N1365);
and AND3 (N5474, N5473, N4853, N4759);
and AND3 (N5475, N5463, N4350, N3157);
and AND2 (N5476, N5470, N472);
xor XOR2 (N5477, N5472, N4690);
buf BUF1 (N5478, N5474);
or OR4 (N5479, N5466, N2569, N4178, N4112);
buf BUF1 (N5480, N5469);
or OR2 (N5481, N5475, N3583);
and AND2 (N5482, N5481, N379);
or OR3 (N5483, N5462, N4527, N2972);
and AND2 (N5484, N5477, N108);
or OR2 (N5485, N5482, N3553);
nor NOR3 (N5486, N5476, N5271, N3279);
and AND3 (N5487, N5467, N5097, N5448);
or OR2 (N5488, N5471, N4355);
nand NAND2 (N5489, N5486, N690);
or OR3 (N5490, N5488, N5215, N4289);
or OR4 (N5491, N5478, N1930, N745, N1710);
xor XOR2 (N5492, N5491, N4015);
xor XOR2 (N5493, N5490, N4296);
and AND4 (N5494, N5479, N3158, N1858, N3109);
buf BUF1 (N5495, N5489);
nand NAND4 (N5496, N5492, N3297, N869, N4788);
nand NAND2 (N5497, N5485, N4651);
not NOT1 (N5498, N5496);
or OR4 (N5499, N5484, N5364, N2047, N723);
nand NAND3 (N5500, N5493, N3866, N1025);
or OR3 (N5501, N5454, N2616, N2679);
and AND4 (N5502, N5500, N1819, N5308, N50);
not NOT1 (N5503, N5502);
or OR2 (N5504, N5480, N5192);
nor NOR4 (N5505, N5494, N1193, N1167, N3052);
or OR4 (N5506, N5501, N4139, N1352, N714);
xor XOR2 (N5507, N5504, N2374);
and AND3 (N5508, N5498, N4783, N3826);
not NOT1 (N5509, N5487);
not NOT1 (N5510, N5507);
nor NOR3 (N5511, N5499, N4907, N1338);
buf BUF1 (N5512, N5508);
xor XOR2 (N5513, N5497, N3542);
or OR3 (N5514, N5510, N1400, N975);
nor NOR3 (N5515, N5511, N1422, N1525);
not NOT1 (N5516, N5512);
nand NAND2 (N5517, N5483, N2961);
nand NAND3 (N5518, N5514, N3872, N3485);
or OR2 (N5519, N5505, N4874);
buf BUF1 (N5520, N5519);
not NOT1 (N5521, N5513);
xor XOR2 (N5522, N5520, N2446);
xor XOR2 (N5523, N5517, N5071);
and AND2 (N5524, N5509, N2596);
nor NOR4 (N5525, N5522, N1824, N4085, N3993);
or OR2 (N5526, N5518, N3537);
buf BUF1 (N5527, N5515);
or OR4 (N5528, N5503, N3772, N1183, N4149);
buf BUF1 (N5529, N5495);
or OR3 (N5530, N5526, N2339, N5420);
nor NOR2 (N5531, N5524, N1080);
not NOT1 (N5532, N5523);
buf BUF1 (N5533, N5525);
nand NAND2 (N5534, N5531, N4885);
xor XOR2 (N5535, N5506, N4360);
not NOT1 (N5536, N5535);
nand NAND2 (N5537, N5536, N3228);
nor NOR4 (N5538, N5521, N3196, N2196, N4987);
nand NAND3 (N5539, N5533, N281, N4743);
not NOT1 (N5540, N5532);
and AND4 (N5541, N5527, N5160, N2608, N5291);
nor NOR2 (N5542, N5530, N3047);
nor NOR3 (N5543, N5534, N3059, N423);
buf BUF1 (N5544, N5538);
nor NOR4 (N5545, N5528, N4769, N344, N3976);
and AND4 (N5546, N5539, N5295, N5481, N1369);
xor XOR2 (N5547, N5541, N5133);
and AND3 (N5548, N5545, N1429, N4743);
nand NAND2 (N5549, N5516, N5244);
buf BUF1 (N5550, N5540);
and AND2 (N5551, N5543, N3675);
not NOT1 (N5552, N5542);
and AND2 (N5553, N5550, N541);
and AND3 (N5554, N5549, N3030, N5247);
xor XOR2 (N5555, N5546, N2144);
or OR4 (N5556, N5552, N3870, N1313, N1449);
or OR2 (N5557, N5537, N3579);
xor XOR2 (N5558, N5554, N2345);
or OR3 (N5559, N5555, N1972, N2737);
and AND4 (N5560, N5547, N4096, N2178, N684);
nand NAND3 (N5561, N5558, N1587, N2736);
buf BUF1 (N5562, N5557);
xor XOR2 (N5563, N5544, N3394);
xor XOR2 (N5564, N5556, N2179);
not NOT1 (N5565, N5560);
or OR4 (N5566, N5551, N720, N1116, N1029);
xor XOR2 (N5567, N5563, N2074);
not NOT1 (N5568, N5553);
nand NAND2 (N5569, N5566, N1577);
and AND2 (N5570, N5561, N665);
and AND2 (N5571, N5567, N4192);
nor NOR4 (N5572, N5564, N2076, N3437, N3419);
or OR3 (N5573, N5569, N5055, N3948);
nor NOR3 (N5574, N5562, N1978, N5212);
and AND4 (N5575, N5574, N1039, N4835, N2665);
nand NAND2 (N5576, N5571, N1898);
not NOT1 (N5577, N5570);
buf BUF1 (N5578, N5573);
nor NOR2 (N5579, N5572, N5537);
nor NOR4 (N5580, N5529, N5057, N654, N3179);
and AND2 (N5581, N5578, N5413);
nand NAND2 (N5582, N5565, N1113);
buf BUF1 (N5583, N5581);
nor NOR2 (N5584, N5548, N3897);
and AND2 (N5585, N5577, N4735);
or OR4 (N5586, N5576, N4758, N4485, N834);
and AND4 (N5587, N5559, N4205, N719, N1946);
nor NOR4 (N5588, N5587, N1783, N148, N3450);
or OR2 (N5589, N5583, N2131);
buf BUF1 (N5590, N5584);
xor XOR2 (N5591, N5575, N2493);
nand NAND4 (N5592, N5585, N2073, N4151, N2978);
nor NOR2 (N5593, N5568, N3678);
not NOT1 (N5594, N5582);
nor NOR2 (N5595, N5589, N3031);
not NOT1 (N5596, N5594);
or OR3 (N5597, N5591, N3443, N5022);
buf BUF1 (N5598, N5586);
and AND2 (N5599, N5598, N3822);
nand NAND2 (N5600, N5588, N3383);
buf BUF1 (N5601, N5596);
xor XOR2 (N5602, N5600, N4256);
not NOT1 (N5603, N5601);
buf BUF1 (N5604, N5592);
buf BUF1 (N5605, N5579);
buf BUF1 (N5606, N5597);
xor XOR2 (N5607, N5580, N340);
xor XOR2 (N5608, N5604, N2946);
not NOT1 (N5609, N5602);
nor NOR4 (N5610, N5603, N2419, N244, N3061);
or OR3 (N5611, N5595, N4739, N2164);
nand NAND4 (N5612, N5605, N1761, N380, N870);
nor NOR4 (N5613, N5590, N973, N1574, N269);
buf BUF1 (N5614, N5612);
buf BUF1 (N5615, N5611);
nand NAND4 (N5616, N5613, N5546, N4937, N1232);
buf BUF1 (N5617, N5608);
xor XOR2 (N5618, N5610, N5365);
nand NAND4 (N5619, N5617, N576, N2833, N4956);
buf BUF1 (N5620, N5619);
not NOT1 (N5621, N5606);
buf BUF1 (N5622, N5607);
xor XOR2 (N5623, N5609, N4002);
buf BUF1 (N5624, N5614);
or OR4 (N5625, N5621, N4352, N2444, N2934);
nor NOR3 (N5626, N5620, N1363, N156);
buf BUF1 (N5627, N5615);
or OR4 (N5628, N5616, N3231, N3158, N319);
xor XOR2 (N5629, N5599, N2040);
not NOT1 (N5630, N5629);
xor XOR2 (N5631, N5624, N1759);
and AND3 (N5632, N5626, N2948, N2755);
xor XOR2 (N5633, N5632, N4018);
or OR4 (N5634, N5630, N4949, N1549, N2499);
nand NAND3 (N5635, N5622, N120, N1178);
xor XOR2 (N5636, N5627, N2664);
buf BUF1 (N5637, N5593);
or OR2 (N5638, N5635, N1228);
nor NOR3 (N5639, N5625, N5347, N2513);
nor NOR4 (N5640, N5634, N2794, N4661, N2745);
xor XOR2 (N5641, N5639, N4283);
buf BUF1 (N5642, N5641);
nor NOR3 (N5643, N5631, N4194, N1035);
nor NOR4 (N5644, N5636, N4120, N4640, N4867);
not NOT1 (N5645, N5633);
not NOT1 (N5646, N5638);
nand NAND4 (N5647, N5640, N3297, N5103, N502);
not NOT1 (N5648, N5643);
not NOT1 (N5649, N5647);
nand NAND4 (N5650, N5646, N610, N5059, N3593);
not NOT1 (N5651, N5645);
xor XOR2 (N5652, N5628, N1478);
xor XOR2 (N5653, N5652, N728);
buf BUF1 (N5654, N5653);
and AND3 (N5655, N5642, N1669, N2952);
nand NAND2 (N5656, N5651, N5215);
and AND2 (N5657, N5618, N2252);
buf BUF1 (N5658, N5644);
xor XOR2 (N5659, N5623, N3078);
not NOT1 (N5660, N5657);
nand NAND4 (N5661, N5648, N4030, N1224, N5539);
and AND3 (N5662, N5656, N4928, N4046);
xor XOR2 (N5663, N5662, N1149);
not NOT1 (N5664, N5655);
buf BUF1 (N5665, N5664);
xor XOR2 (N5666, N5665, N4882);
xor XOR2 (N5667, N5650, N5290);
not NOT1 (N5668, N5661);
not NOT1 (N5669, N5658);
nand NAND4 (N5670, N5660, N1804, N3923, N5192);
buf BUF1 (N5671, N5668);
nor NOR2 (N5672, N5663, N3307);
nand NAND4 (N5673, N5670, N5194, N3714, N5204);
buf BUF1 (N5674, N5666);
not NOT1 (N5675, N5673);
not NOT1 (N5676, N5672);
nor NOR2 (N5677, N5671, N5657);
nand NAND2 (N5678, N5675, N4650);
or OR3 (N5679, N5637, N2992, N4834);
not NOT1 (N5680, N5677);
and AND4 (N5681, N5659, N2500, N710, N501);
nand NAND2 (N5682, N5667, N4430);
and AND4 (N5683, N5654, N3615, N3996, N2811);
not NOT1 (N5684, N5674);
buf BUF1 (N5685, N5669);
not NOT1 (N5686, N5678);
buf BUF1 (N5687, N5676);
not NOT1 (N5688, N5680);
and AND3 (N5689, N5688, N3424, N1291);
nand NAND4 (N5690, N5681, N3754, N322, N208);
or OR3 (N5691, N5679, N5506, N4977);
or OR4 (N5692, N5689, N631, N378, N2867);
xor XOR2 (N5693, N5691, N295);
nand NAND4 (N5694, N5692, N3803, N3907, N2773);
nor NOR3 (N5695, N5684, N3643, N2670);
nor NOR3 (N5696, N5694, N600, N4419);
buf BUF1 (N5697, N5685);
and AND2 (N5698, N5687, N5551);
not NOT1 (N5699, N5696);
xor XOR2 (N5700, N5699, N2501);
nor NOR3 (N5701, N5683, N4928, N2873);
nor NOR3 (N5702, N5690, N1484, N4199);
and AND4 (N5703, N5695, N2782, N4599, N3178);
or OR4 (N5704, N5649, N3728, N1467, N1419);
and AND3 (N5705, N5701, N384, N199);
or OR4 (N5706, N5702, N1904, N3755, N4956);
nand NAND2 (N5707, N5686, N3941);
buf BUF1 (N5708, N5706);
and AND2 (N5709, N5707, N3633);
and AND3 (N5710, N5697, N4247, N939);
or OR2 (N5711, N5703, N5074);
not NOT1 (N5712, N5710);
not NOT1 (N5713, N5693);
and AND4 (N5714, N5709, N3861, N2211, N4408);
xor XOR2 (N5715, N5712, N403);
or OR4 (N5716, N5700, N762, N2738, N4230);
nand NAND2 (N5717, N5704, N5028);
xor XOR2 (N5718, N5708, N5261);
nand NAND4 (N5719, N5715, N1384, N5307, N1777);
buf BUF1 (N5720, N5698);
or OR3 (N5721, N5717, N4679, N2655);
xor XOR2 (N5722, N5713, N3814);
nand NAND3 (N5723, N5722, N4490, N4984);
nor NOR4 (N5724, N5718, N3651, N5074, N3284);
nor NOR4 (N5725, N5724, N726, N4464, N1688);
or OR2 (N5726, N5682, N1698);
or OR4 (N5727, N5726, N421, N5199, N88);
nand NAND3 (N5728, N5711, N2626, N4261);
or OR3 (N5729, N5721, N1725, N1469);
or OR2 (N5730, N5714, N2093);
or OR4 (N5731, N5729, N2202, N4463, N1911);
and AND2 (N5732, N5719, N1645);
nor NOR4 (N5733, N5720, N5649, N3419, N3823);
and AND2 (N5734, N5730, N2967);
xor XOR2 (N5735, N5733, N4661);
xor XOR2 (N5736, N5732, N2409);
xor XOR2 (N5737, N5705, N2415);
nand NAND3 (N5738, N5728, N4860, N3778);
nor NOR3 (N5739, N5734, N1650, N5374);
or OR4 (N5740, N5731, N5068, N835, N4995);
nand NAND4 (N5741, N5725, N2236, N3522, N4668);
nor NOR2 (N5742, N5723, N3695);
and AND4 (N5743, N5736, N4265, N78, N1734);
or OR2 (N5744, N5737, N2589);
buf BUF1 (N5745, N5739);
nor NOR2 (N5746, N5744, N3172);
nand NAND3 (N5747, N5746, N4903, N4569);
or OR4 (N5748, N5716, N5218, N3579, N1271);
nor NOR4 (N5749, N5741, N2951, N2889, N244);
buf BUF1 (N5750, N5742);
or OR2 (N5751, N5750, N3123);
nor NOR4 (N5752, N5748, N1539, N5550, N4023);
and AND2 (N5753, N5749, N989);
buf BUF1 (N5754, N5753);
nor NOR4 (N5755, N5738, N2019, N2017, N830);
not NOT1 (N5756, N5755);
not NOT1 (N5757, N5745);
nand NAND2 (N5758, N5740, N1538);
buf BUF1 (N5759, N5735);
not NOT1 (N5760, N5751);
buf BUF1 (N5761, N5754);
xor XOR2 (N5762, N5743, N5418);
and AND3 (N5763, N5752, N1059, N4888);
xor XOR2 (N5764, N5758, N1801);
and AND2 (N5765, N5761, N1245);
nor NOR2 (N5766, N5756, N2609);
xor XOR2 (N5767, N5757, N4552);
xor XOR2 (N5768, N5767, N2870);
not NOT1 (N5769, N5768);
xor XOR2 (N5770, N5766, N5233);
and AND4 (N5771, N5760, N4531, N4737, N1255);
not NOT1 (N5772, N5769);
buf BUF1 (N5773, N5770);
nand NAND3 (N5774, N5747, N2444, N1337);
nand NAND2 (N5775, N5765, N1576);
not NOT1 (N5776, N5773);
or OR3 (N5777, N5759, N5749, N2312);
or OR3 (N5778, N5727, N5760, N322);
buf BUF1 (N5779, N5776);
and AND3 (N5780, N5779, N169, N1704);
buf BUF1 (N5781, N5774);
or OR2 (N5782, N5781, N1744);
not NOT1 (N5783, N5764);
buf BUF1 (N5784, N5777);
not NOT1 (N5785, N5771);
or OR4 (N5786, N5763, N4526, N1539, N3433);
buf BUF1 (N5787, N5783);
xor XOR2 (N5788, N5784, N1547);
nand NAND2 (N5789, N5785, N4922);
buf BUF1 (N5790, N5772);
nand NAND4 (N5791, N5775, N184, N5735, N2051);
nand NAND4 (N5792, N5791, N4340, N3823, N498);
xor XOR2 (N5793, N5782, N1004);
not NOT1 (N5794, N5787);
nand NAND4 (N5795, N5793, N3109, N5643, N4762);
nand NAND2 (N5796, N5788, N1601);
and AND4 (N5797, N5789, N5515, N3487, N3455);
nor NOR2 (N5798, N5794, N4528);
xor XOR2 (N5799, N5786, N5434);
and AND4 (N5800, N5762, N4571, N2295, N5128);
buf BUF1 (N5801, N5797);
or OR2 (N5802, N5801, N5716);
xor XOR2 (N5803, N5796, N1535);
xor XOR2 (N5804, N5778, N4289);
nor NOR4 (N5805, N5790, N3953, N3767, N954);
xor XOR2 (N5806, N5798, N3492);
and AND4 (N5807, N5802, N4450, N1021, N2494);
not NOT1 (N5808, N5806);
buf BUF1 (N5809, N5803);
not NOT1 (N5810, N5800);
nand NAND2 (N5811, N5780, N2583);
and AND2 (N5812, N5807, N1832);
and AND2 (N5813, N5811, N2345);
xor XOR2 (N5814, N5809, N4733);
or OR3 (N5815, N5813, N3060, N2520);
buf BUF1 (N5816, N5815);
and AND3 (N5817, N5799, N4507, N4442);
not NOT1 (N5818, N5810);
nor NOR2 (N5819, N5805, N2852);
xor XOR2 (N5820, N5795, N1076);
or OR4 (N5821, N5816, N693, N5626, N1812);
xor XOR2 (N5822, N5814, N2123);
not NOT1 (N5823, N5821);
not NOT1 (N5824, N5818);
nand NAND3 (N5825, N5812, N4645, N4346);
nand NAND2 (N5826, N5824, N5194);
not NOT1 (N5827, N5822);
buf BUF1 (N5828, N5820);
or OR3 (N5829, N5826, N2356, N2905);
or OR4 (N5830, N5827, N5572, N2135, N2071);
or OR3 (N5831, N5819, N1970, N1015);
and AND4 (N5832, N5825, N2059, N4982, N4945);
and AND2 (N5833, N5817, N647);
buf BUF1 (N5834, N5831);
or OR2 (N5835, N5834, N5706);
and AND3 (N5836, N5792, N4019, N1421);
not NOT1 (N5837, N5808);
nand NAND4 (N5838, N5823, N5102, N2988, N5259);
not NOT1 (N5839, N5832);
not NOT1 (N5840, N5804);
xor XOR2 (N5841, N5839, N4832);
buf BUF1 (N5842, N5837);
buf BUF1 (N5843, N5840);
nand NAND4 (N5844, N5828, N5603, N4561, N392);
and AND4 (N5845, N5842, N4127, N2640, N2674);
xor XOR2 (N5846, N5838, N2751);
xor XOR2 (N5847, N5829, N3089);
xor XOR2 (N5848, N5841, N1219);
not NOT1 (N5849, N5844);
buf BUF1 (N5850, N5848);
xor XOR2 (N5851, N5845, N1088);
not NOT1 (N5852, N5833);
nor NOR4 (N5853, N5852, N1756, N174, N3500);
or OR4 (N5854, N5830, N3901, N5643, N3029);
nor NOR4 (N5855, N5854, N4957, N4531, N331);
not NOT1 (N5856, N5846);
buf BUF1 (N5857, N5851);
nand NAND4 (N5858, N5847, N311, N4839, N3069);
buf BUF1 (N5859, N5843);
nand NAND4 (N5860, N5857, N4056, N4180, N3333);
and AND3 (N5861, N5855, N4967, N4382);
or OR3 (N5862, N5861, N3803, N5176);
nand NAND2 (N5863, N5858, N5049);
or OR2 (N5864, N5862, N215);
or OR4 (N5865, N5856, N4661, N3926, N4654);
not NOT1 (N5866, N5850);
nor NOR3 (N5867, N5853, N147, N1766);
or OR4 (N5868, N5860, N2641, N3840, N3458);
buf BUF1 (N5869, N5866);
nand NAND3 (N5870, N5865, N1093, N1800);
nor NOR4 (N5871, N5859, N2946, N1980, N4661);
and AND3 (N5872, N5835, N1567, N4453);
xor XOR2 (N5873, N5867, N1846);
xor XOR2 (N5874, N5870, N2870);
or OR4 (N5875, N5869, N2216, N3470, N1799);
and AND2 (N5876, N5836, N3084);
buf BUF1 (N5877, N5849);
xor XOR2 (N5878, N5872, N17);
buf BUF1 (N5879, N5878);
not NOT1 (N5880, N5868);
or OR2 (N5881, N5875, N1750);
xor XOR2 (N5882, N5880, N2121);
nand NAND4 (N5883, N5873, N385, N5021, N1109);
and AND4 (N5884, N5864, N3694, N1063, N1395);
xor XOR2 (N5885, N5877, N1581);
not NOT1 (N5886, N5871);
xor XOR2 (N5887, N5885, N5802);
nand NAND2 (N5888, N5886, N4646);
buf BUF1 (N5889, N5876);
and AND3 (N5890, N5879, N4538, N3812);
and AND2 (N5891, N5888, N5220);
nor NOR4 (N5892, N5883, N137, N2132, N3635);
xor XOR2 (N5893, N5887, N2697);
buf BUF1 (N5894, N5884);
nand NAND4 (N5895, N5874, N4508, N4358, N2090);
and AND4 (N5896, N5890, N3820, N1243, N2172);
nor NOR3 (N5897, N5891, N41, N590);
buf BUF1 (N5898, N5881);
buf BUF1 (N5899, N5898);
not NOT1 (N5900, N5892);
xor XOR2 (N5901, N5863, N5399);
buf BUF1 (N5902, N5882);
not NOT1 (N5903, N5897);
or OR2 (N5904, N5899, N5234);
and AND4 (N5905, N5900, N2778, N1463, N1559);
xor XOR2 (N5906, N5901, N5901);
or OR4 (N5907, N5903, N2975, N3581, N4076);
nor NOR2 (N5908, N5907, N5300);
and AND4 (N5909, N5906, N5178, N736, N5707);
nor NOR2 (N5910, N5905, N3670);
xor XOR2 (N5911, N5908, N952);
buf BUF1 (N5912, N5902);
or OR2 (N5913, N5912, N3005);
xor XOR2 (N5914, N5910, N2494);
xor XOR2 (N5915, N5896, N4243);
and AND4 (N5916, N5904, N4505, N288, N5715);
and AND4 (N5917, N5895, N242, N2234, N4973);
nand NAND4 (N5918, N5909, N1159, N1577, N1219);
nand NAND3 (N5919, N5913, N5740, N1404);
nand NAND2 (N5920, N5889, N1752);
and AND4 (N5921, N5917, N5480, N5393, N5907);
nand NAND3 (N5922, N5916, N1134, N1008);
and AND3 (N5923, N5915, N2217, N5564);
nor NOR4 (N5924, N5894, N3110, N5683, N3108);
nand NAND4 (N5925, N5911, N4445, N4702, N233);
not NOT1 (N5926, N5920);
buf BUF1 (N5927, N5922);
or OR3 (N5928, N5921, N3876, N4591);
and AND2 (N5929, N5918, N5170);
nand NAND4 (N5930, N5926, N2234, N4727, N264);
or OR3 (N5931, N5919, N3132, N4881);
nand NAND2 (N5932, N5925, N4564);
not NOT1 (N5933, N5929);
not NOT1 (N5934, N5932);
xor XOR2 (N5935, N5928, N4049);
nand NAND4 (N5936, N5935, N2370, N2161, N1539);
and AND4 (N5937, N5930, N5065, N3061, N2411);
nand NAND3 (N5938, N5936, N4000, N1341);
xor XOR2 (N5939, N5933, N5308);
or OR2 (N5940, N5931, N534);
and AND2 (N5941, N5924, N4681);
nand NAND4 (N5942, N5914, N5462, N322, N1637);
buf BUF1 (N5943, N5923);
buf BUF1 (N5944, N5927);
xor XOR2 (N5945, N5939, N5299);
or OR4 (N5946, N5934, N3157, N5064, N2595);
not NOT1 (N5947, N5938);
nor NOR4 (N5948, N5941, N2178, N5513, N4948);
nor NOR3 (N5949, N5942, N404, N289);
and AND4 (N5950, N5945, N1769, N5218, N3525);
nand NAND3 (N5951, N5944, N5452, N1429);
nand NAND4 (N5952, N5937, N1547, N2322, N3395);
xor XOR2 (N5953, N5943, N5474);
or OR2 (N5954, N5951, N4517);
and AND4 (N5955, N5954, N986, N1525, N5890);
or OR3 (N5956, N5946, N395, N4410);
not NOT1 (N5957, N5947);
nand NAND4 (N5958, N5953, N1745, N284, N745);
or OR3 (N5959, N5949, N931, N2023);
and AND3 (N5960, N5956, N5532, N2181);
nor NOR4 (N5961, N5893, N2174, N3379, N5650);
and AND3 (N5962, N5960, N4428, N323);
and AND4 (N5963, N5955, N4217, N1847, N1588);
not NOT1 (N5964, N5958);
and AND3 (N5965, N5962, N2041, N4686);
or OR4 (N5966, N5964, N5785, N5751, N4199);
buf BUF1 (N5967, N5965);
and AND2 (N5968, N5961, N3305);
or OR3 (N5969, N5950, N514, N172);
nand NAND3 (N5970, N5959, N4191, N5077);
not NOT1 (N5971, N5966);
nand NAND2 (N5972, N5969, N1926);
not NOT1 (N5973, N5970);
or OR3 (N5974, N5963, N535, N4126);
not NOT1 (N5975, N5967);
nand NAND3 (N5976, N5968, N5507, N3356);
and AND3 (N5977, N5948, N5667, N3328);
and AND4 (N5978, N5972, N3765, N2504, N3832);
or OR3 (N5979, N5940, N5108, N4481);
not NOT1 (N5980, N5979);
or OR3 (N5981, N5975, N3736, N3238);
not NOT1 (N5982, N5957);
nor NOR2 (N5983, N5976, N5544);
buf BUF1 (N5984, N5983);
buf BUF1 (N5985, N5977);
nor NOR2 (N5986, N5984, N1008);
not NOT1 (N5987, N5978);
not NOT1 (N5988, N5986);
or OR3 (N5989, N5981, N3387, N2653);
nand NAND2 (N5990, N5973, N1730);
xor XOR2 (N5991, N5985, N4732);
and AND4 (N5992, N5974, N2810, N5437, N4906);
nor NOR2 (N5993, N5989, N5600);
or OR2 (N5994, N5980, N236);
not NOT1 (N5995, N5994);
and AND3 (N5996, N5971, N2067, N2571);
or OR2 (N5997, N5993, N5526);
or OR4 (N5998, N5995, N2389, N3685, N4782);
or OR4 (N5999, N5998, N1274, N5632, N961);
nand NAND3 (N6000, N5990, N1895, N1953);
and AND4 (N6001, N5982, N2272, N2553, N1225);
or OR4 (N6002, N6000, N5505, N2272, N2292);
or OR4 (N6003, N6001, N998, N5207, N842);
nor NOR3 (N6004, N5988, N5147, N2037);
buf BUF1 (N6005, N6003);
nand NAND3 (N6006, N5999, N406, N5833);
or OR3 (N6007, N6004, N5321, N1251);
not NOT1 (N6008, N6002);
nor NOR4 (N6009, N5991, N5670, N2554, N4489);
or OR2 (N6010, N6008, N1980);
nand NAND3 (N6011, N6007, N1597, N1370);
nand NAND3 (N6012, N5987, N4245, N4279);
xor XOR2 (N6013, N5997, N5630);
and AND2 (N6014, N6013, N5704);
nand NAND4 (N6015, N6005, N2321, N3888, N5004);
and AND3 (N6016, N5952, N2660, N1473);
or OR3 (N6017, N6009, N4914, N4893);
not NOT1 (N6018, N6012);
nand NAND2 (N6019, N6017, N2734);
xor XOR2 (N6020, N6015, N1830);
nand NAND2 (N6021, N6006, N1674);
xor XOR2 (N6022, N6018, N3973);
nor NOR4 (N6023, N6011, N5330, N3400, N2923);
and AND2 (N6024, N5996, N4804);
not NOT1 (N6025, N6019);
nor NOR3 (N6026, N5992, N4060, N636);
nand NAND4 (N6027, N6014, N4168, N1212, N176);
xor XOR2 (N6028, N6010, N5282);
nand NAND3 (N6029, N6020, N5324, N1605);
and AND3 (N6030, N6016, N4, N5630);
not NOT1 (N6031, N6028);
or OR4 (N6032, N6027, N1109, N1235, N1718);
nand NAND4 (N6033, N6026, N6008, N812, N4460);
not NOT1 (N6034, N6023);
or OR3 (N6035, N6031, N790, N1201);
buf BUF1 (N6036, N6024);
or OR4 (N6037, N6034, N418, N1320, N4596);
xor XOR2 (N6038, N6021, N4742);
nor NOR4 (N6039, N6032, N5271, N6023, N5594);
xor XOR2 (N6040, N6022, N5040);
not NOT1 (N6041, N6040);
nor NOR3 (N6042, N6033, N5398, N4078);
nor NOR2 (N6043, N6041, N3120);
nor NOR3 (N6044, N6029, N5036, N2044);
buf BUF1 (N6045, N6043);
and AND3 (N6046, N6044, N176, N2511);
nand NAND4 (N6047, N6038, N5888, N5961, N2597);
or OR2 (N6048, N6042, N2918);
and AND3 (N6049, N6039, N782, N4509);
nand NAND4 (N6050, N6048, N4259, N3579, N5308);
xor XOR2 (N6051, N6036, N596);
and AND3 (N6052, N6049, N2801, N2844);
buf BUF1 (N6053, N6046);
buf BUF1 (N6054, N6030);
xor XOR2 (N6055, N6052, N1988);
not NOT1 (N6056, N6054);
and AND2 (N6057, N6037, N4556);
xor XOR2 (N6058, N6057, N5628);
xor XOR2 (N6059, N6055, N2473);
nand NAND2 (N6060, N6051, N1259);
and AND4 (N6061, N6047, N4865, N1618, N5178);
or OR2 (N6062, N6060, N5815);
or OR3 (N6063, N6045, N2022, N1608);
nand NAND4 (N6064, N6058, N3040, N4913, N996);
nand NAND3 (N6065, N6061, N954, N4380);
nor NOR2 (N6066, N6064, N5013);
xor XOR2 (N6067, N6053, N3155);
nand NAND2 (N6068, N6067, N73);
buf BUF1 (N6069, N6059);
not NOT1 (N6070, N6069);
and AND4 (N6071, N6056, N1211, N3339, N724);
nand NAND2 (N6072, N6068, N1074);
not NOT1 (N6073, N6066);
or OR2 (N6074, N6050, N4254);
xor XOR2 (N6075, N6065, N1566);
and AND4 (N6076, N6072, N1183, N4106, N4276);
nor NOR2 (N6077, N6062, N563);
buf BUF1 (N6078, N6076);
nand NAND3 (N6079, N6070, N2936, N3226);
or OR3 (N6080, N6073, N1032, N2018);
nor NOR2 (N6081, N6063, N2407);
and AND3 (N6082, N6071, N4628, N5107);
or OR2 (N6083, N6079, N4544);
and AND4 (N6084, N6025, N3586, N5168, N1681);
buf BUF1 (N6085, N6077);
buf BUF1 (N6086, N6035);
nor NOR4 (N6087, N6083, N5586, N731, N1758);
nor NOR3 (N6088, N6081, N3786, N4938);
nand NAND4 (N6089, N6080, N1870, N3927, N5239);
xor XOR2 (N6090, N6085, N1402);
buf BUF1 (N6091, N6086);
xor XOR2 (N6092, N6090, N3103);
nor NOR3 (N6093, N6074, N2059, N3770);
buf BUF1 (N6094, N6092);
nor NOR3 (N6095, N6084, N2047, N2683);
nand NAND4 (N6096, N6087, N2663, N4589, N2516);
not NOT1 (N6097, N6091);
nor NOR4 (N6098, N6075, N1804, N2200, N1178);
nor NOR3 (N6099, N6089, N5845, N367);
buf BUF1 (N6100, N6099);
nor NOR3 (N6101, N6098, N412, N4649);
and AND4 (N6102, N6101, N2401, N4366, N3153);
and AND4 (N6103, N6102, N1240, N4053, N2982);
buf BUF1 (N6104, N6088);
and AND4 (N6105, N6103, N5758, N3541, N3270);
nand NAND4 (N6106, N6100, N5326, N3029, N4724);
buf BUF1 (N6107, N6106);
nand NAND2 (N6108, N6105, N2321);
nor NOR2 (N6109, N6078, N5879);
buf BUF1 (N6110, N6093);
and AND2 (N6111, N6104, N5723);
or OR3 (N6112, N6111, N1605, N4348);
or OR2 (N6113, N6096, N3567);
buf BUF1 (N6114, N6109);
and AND3 (N6115, N6114, N5877, N2373);
nand NAND2 (N6116, N6094, N5057);
not NOT1 (N6117, N6113);
not NOT1 (N6118, N6117);
and AND3 (N6119, N6095, N4567, N3826);
xor XOR2 (N6120, N6115, N5807);
nand NAND2 (N6121, N6116, N2900);
nor NOR3 (N6122, N6119, N2204, N5958);
nor NOR4 (N6123, N6082, N471, N3499, N1901);
or OR4 (N6124, N6121, N5715, N1966, N3422);
not NOT1 (N6125, N6124);
buf BUF1 (N6126, N6097);
buf BUF1 (N6127, N6107);
buf BUF1 (N6128, N6127);
or OR2 (N6129, N6110, N3152);
xor XOR2 (N6130, N6128, N5816);
buf BUF1 (N6131, N6126);
or OR4 (N6132, N6131, N3517, N3440, N82);
xor XOR2 (N6133, N6112, N5674);
xor XOR2 (N6134, N6123, N3795);
nand NAND2 (N6135, N6108, N3926);
not NOT1 (N6136, N6134);
buf BUF1 (N6137, N6125);
xor XOR2 (N6138, N6120, N5211);
buf BUF1 (N6139, N6130);
and AND3 (N6140, N6118, N3543, N3806);
nand NAND3 (N6141, N6138, N1416, N688);
xor XOR2 (N6142, N6129, N696);
not NOT1 (N6143, N6136);
or OR3 (N6144, N6142, N525, N2801);
not NOT1 (N6145, N6137);
or OR4 (N6146, N6145, N5593, N5867, N2674);
or OR4 (N6147, N6144, N3734, N1146, N3765);
not NOT1 (N6148, N6147);
xor XOR2 (N6149, N6148, N674);
xor XOR2 (N6150, N6149, N2914);
or OR2 (N6151, N6141, N2383);
xor XOR2 (N6152, N6146, N3851);
nor NOR4 (N6153, N6150, N1904, N818, N4441);
not NOT1 (N6154, N6140);
and AND2 (N6155, N6139, N1260);
nor NOR3 (N6156, N6143, N5969, N2955);
buf BUF1 (N6157, N6153);
or OR4 (N6158, N6155, N1085, N4756, N4712);
nand NAND2 (N6159, N6158, N2316);
buf BUF1 (N6160, N6157);
nand NAND3 (N6161, N6152, N1030, N5211);
and AND2 (N6162, N6133, N1575);
or OR2 (N6163, N6122, N3806);
nor NOR3 (N6164, N6163, N2345, N4295);
and AND2 (N6165, N6164, N5575);
not NOT1 (N6166, N6154);
not NOT1 (N6167, N6156);
nand NAND4 (N6168, N6167, N2378, N3315, N540);
nor NOR3 (N6169, N6132, N5444, N5291);
buf BUF1 (N6170, N6169);
nor NOR2 (N6171, N6165, N5931);
nand NAND3 (N6172, N6168, N3331, N4171);
nand NAND4 (N6173, N6166, N5343, N4345, N3360);
nor NOR4 (N6174, N6135, N4421, N1149, N3719);
nor NOR4 (N6175, N6161, N3430, N4624, N2344);
buf BUF1 (N6176, N6172);
not NOT1 (N6177, N6176);
xor XOR2 (N6178, N6170, N5416);
not NOT1 (N6179, N6177);
buf BUF1 (N6180, N6179);
nor NOR2 (N6181, N6174, N3673);
or OR2 (N6182, N6151, N4859);
buf BUF1 (N6183, N6173);
nand NAND2 (N6184, N6181, N1280);
xor XOR2 (N6185, N6184, N1978);
nor NOR4 (N6186, N6182, N1032, N4069, N2626);
not NOT1 (N6187, N6183);
buf BUF1 (N6188, N6175);
not NOT1 (N6189, N6159);
and AND4 (N6190, N6189, N1319, N2877, N3871);
nor NOR2 (N6191, N6160, N2999);
nand NAND3 (N6192, N6187, N5746, N1947);
buf BUF1 (N6193, N6162);
buf BUF1 (N6194, N6191);
not NOT1 (N6195, N6192);
xor XOR2 (N6196, N6190, N1639);
or OR2 (N6197, N6171, N3274);
xor XOR2 (N6198, N6196, N4723);
not NOT1 (N6199, N6194);
nor NOR2 (N6200, N6188, N54);
buf BUF1 (N6201, N6198);
nor NOR3 (N6202, N6193, N5934, N4068);
and AND3 (N6203, N6195, N5186, N1875);
buf BUF1 (N6204, N6200);
nor NOR4 (N6205, N6202, N2028, N124, N3122);
nand NAND4 (N6206, N6186, N5922, N5390, N5862);
or OR3 (N6207, N6206, N4768, N4733);
or OR2 (N6208, N6180, N3510);
not NOT1 (N6209, N6199);
buf BUF1 (N6210, N6178);
not NOT1 (N6211, N6205);
not NOT1 (N6212, N6201);
not NOT1 (N6213, N6185);
buf BUF1 (N6214, N6211);
or OR4 (N6215, N6214, N1072, N2760, N5392);
not NOT1 (N6216, N6210);
xor XOR2 (N6217, N6203, N1064);
xor XOR2 (N6218, N6215, N3413);
nor NOR2 (N6219, N6197, N5915);
not NOT1 (N6220, N6216);
nor NOR3 (N6221, N6217, N4664, N2931);
or OR3 (N6222, N6209, N5745, N6);
not NOT1 (N6223, N6219);
and AND2 (N6224, N6218, N1023);
and AND3 (N6225, N6224, N109, N2204);
and AND3 (N6226, N6225, N2447, N6099);
nand NAND4 (N6227, N6220, N2298, N2299, N6159);
nand NAND2 (N6228, N6204, N117);
buf BUF1 (N6229, N6221);
nand NAND3 (N6230, N6208, N4148, N1471);
not NOT1 (N6231, N6223);
buf BUF1 (N6232, N6222);
and AND2 (N6233, N6227, N5989);
not NOT1 (N6234, N6230);
xor XOR2 (N6235, N6207, N3864);
or OR4 (N6236, N6231, N986, N1390, N2339);
nor NOR2 (N6237, N6228, N1862);
buf BUF1 (N6238, N6213);
nand NAND4 (N6239, N6234, N943, N3763, N3100);
nand NAND4 (N6240, N6212, N3499, N3863, N2981);
buf BUF1 (N6241, N6226);
not NOT1 (N6242, N6229);
not NOT1 (N6243, N6237);
nor NOR2 (N6244, N6232, N5914);
or OR4 (N6245, N6238, N4819, N5806, N4704);
buf BUF1 (N6246, N6245);
not NOT1 (N6247, N6239);
and AND3 (N6248, N6241, N6053, N5054);
and AND4 (N6249, N6240, N5051, N14, N320);
or OR3 (N6250, N6244, N5314, N91);
xor XOR2 (N6251, N6250, N3703);
buf BUF1 (N6252, N6243);
not NOT1 (N6253, N6235);
not NOT1 (N6254, N6242);
nor NOR3 (N6255, N6251, N3358, N2385);
and AND4 (N6256, N6248, N5769, N3119, N3574);
buf BUF1 (N6257, N6256);
and AND3 (N6258, N6257, N3918, N2027);
buf BUF1 (N6259, N6236);
nor NOR4 (N6260, N6258, N4787, N2475, N4103);
not NOT1 (N6261, N6249);
buf BUF1 (N6262, N6261);
nand NAND4 (N6263, N6253, N3177, N3096, N5772);
xor XOR2 (N6264, N6254, N3617);
or OR2 (N6265, N6263, N383);
and AND3 (N6266, N6247, N3089, N5879);
not NOT1 (N6267, N6233);
xor XOR2 (N6268, N6262, N2347);
buf BUF1 (N6269, N6266);
xor XOR2 (N6270, N6255, N5494);
not NOT1 (N6271, N6267);
not NOT1 (N6272, N6269);
buf BUF1 (N6273, N6252);
and AND2 (N6274, N6273, N1099);
xor XOR2 (N6275, N6265, N2476);
buf BUF1 (N6276, N6264);
or OR3 (N6277, N6275, N2444, N2514);
nor NOR2 (N6278, N6276, N5921);
not NOT1 (N6279, N6274);
nor NOR3 (N6280, N6268, N4146, N398);
xor XOR2 (N6281, N6259, N2443);
xor XOR2 (N6282, N6281, N2344);
not NOT1 (N6283, N6277);
buf BUF1 (N6284, N6260);
buf BUF1 (N6285, N6284);
xor XOR2 (N6286, N6285, N4426);
buf BUF1 (N6287, N6283);
nand NAND3 (N6288, N6270, N5275, N2028);
not NOT1 (N6289, N6280);
nor NOR3 (N6290, N6271, N3083, N5559);
xor XOR2 (N6291, N6287, N3694);
or OR4 (N6292, N6288, N1850, N2347, N5165);
or OR4 (N6293, N6291, N5035, N1531, N192);
nand NAND4 (N6294, N6272, N2402, N3078, N224);
nor NOR2 (N6295, N6292, N3377);
buf BUF1 (N6296, N6286);
or OR3 (N6297, N6289, N4760, N1246);
not NOT1 (N6298, N6282);
nand NAND3 (N6299, N6293, N2669, N1811);
not NOT1 (N6300, N6299);
nand NAND2 (N6301, N6300, N1175);
buf BUF1 (N6302, N6296);
or OR2 (N6303, N6290, N848);
buf BUF1 (N6304, N6298);
xor XOR2 (N6305, N6246, N2150);
nor NOR3 (N6306, N6305, N5219, N3276);
nor NOR3 (N6307, N6297, N4767, N1045);
and AND3 (N6308, N6304, N3082, N1658);
nor NOR4 (N6309, N6294, N1045, N1387, N4589);
buf BUF1 (N6310, N6309);
nand NAND3 (N6311, N6307, N3524, N3676);
not NOT1 (N6312, N6308);
not NOT1 (N6313, N6279);
not NOT1 (N6314, N6302);
nand NAND2 (N6315, N6314, N2674);
xor XOR2 (N6316, N6312, N1764);
or OR2 (N6317, N6295, N4767);
buf BUF1 (N6318, N6317);
not NOT1 (N6319, N6310);
nand NAND3 (N6320, N6318, N4656, N5746);
nand NAND2 (N6321, N6313, N3865);
not NOT1 (N6322, N6315);
nor NOR2 (N6323, N6278, N4757);
nand NAND2 (N6324, N6301, N3774);
and AND4 (N6325, N6306, N975, N6073, N4773);
and AND2 (N6326, N6311, N838);
xor XOR2 (N6327, N6316, N6052);
and AND4 (N6328, N6323, N739, N5399, N5822);
not NOT1 (N6329, N6324);
and AND2 (N6330, N6319, N2163);
nand NAND2 (N6331, N6325, N1533);
or OR4 (N6332, N6321, N4751, N2172, N254);
buf BUF1 (N6333, N6332);
and AND2 (N6334, N6326, N211);
nand NAND2 (N6335, N6330, N1103);
buf BUF1 (N6336, N6331);
buf BUF1 (N6337, N6335);
and AND3 (N6338, N6333, N1484, N1693);
nor NOR4 (N6339, N6320, N2807, N1263, N4365);
or OR4 (N6340, N6339, N767, N246, N1795);
or OR4 (N6341, N6327, N1550, N2947, N3031);
not NOT1 (N6342, N6340);
nand NAND3 (N6343, N6337, N277, N4709);
or OR4 (N6344, N6334, N2442, N871, N2239);
or OR4 (N6345, N6341, N4591, N3085, N6116);
buf BUF1 (N6346, N6338);
or OR2 (N6347, N6346, N2855);
xor XOR2 (N6348, N6336, N5358);
buf BUF1 (N6349, N6347);
buf BUF1 (N6350, N6342);
xor XOR2 (N6351, N6350, N2781);
or OR4 (N6352, N6345, N1859, N984, N3246);
not NOT1 (N6353, N6351);
not NOT1 (N6354, N6353);
buf BUF1 (N6355, N6344);
buf BUF1 (N6356, N6354);
nor NOR4 (N6357, N6348, N1796, N5477, N3423);
nor NOR2 (N6358, N6349, N2037);
nor NOR2 (N6359, N6356, N390);
xor XOR2 (N6360, N6358, N6125);
and AND2 (N6361, N6303, N4060);
buf BUF1 (N6362, N6361);
not NOT1 (N6363, N6359);
and AND4 (N6364, N6352, N195, N1413, N3579);
buf BUF1 (N6365, N6360);
nand NAND2 (N6366, N6328, N2444);
buf BUF1 (N6367, N6355);
or OR2 (N6368, N6363, N2447);
buf BUF1 (N6369, N6343);
nor NOR2 (N6370, N6362, N2225);
nor NOR3 (N6371, N6368, N4182, N2919);
xor XOR2 (N6372, N6329, N4449);
nand NAND3 (N6373, N6367, N5118, N5309);
buf BUF1 (N6374, N6364);
nor NOR4 (N6375, N6370, N5407, N3518, N6273);
nand NAND2 (N6376, N6375, N6190);
nand NAND3 (N6377, N6365, N5953, N5695);
not NOT1 (N6378, N6371);
or OR2 (N6379, N6373, N1021);
nand NAND4 (N6380, N6366, N3536, N1921, N3129);
xor XOR2 (N6381, N6378, N5898);
buf BUF1 (N6382, N6377);
buf BUF1 (N6383, N6379);
buf BUF1 (N6384, N6376);
xor XOR2 (N6385, N6369, N1888);
and AND2 (N6386, N6384, N3660);
nand NAND4 (N6387, N6385, N3577, N2596, N368);
not NOT1 (N6388, N6372);
not NOT1 (N6389, N6386);
and AND4 (N6390, N6389, N6115, N4356, N4812);
nand NAND2 (N6391, N6357, N396);
xor XOR2 (N6392, N6381, N1455);
nand NAND2 (N6393, N6387, N3534);
buf BUF1 (N6394, N6391);
and AND4 (N6395, N6388, N6069, N3816, N1403);
and AND2 (N6396, N6383, N5461);
and AND2 (N6397, N6390, N1672);
or OR2 (N6398, N6397, N3029);
nand NAND2 (N6399, N6394, N5473);
buf BUF1 (N6400, N6382);
nand NAND4 (N6401, N6395, N258, N409, N5114);
nand NAND3 (N6402, N6392, N2524, N2966);
nor NOR3 (N6403, N6400, N1642, N187);
xor XOR2 (N6404, N6396, N6162);
nor NOR2 (N6405, N6398, N6006);
or OR2 (N6406, N6401, N5480);
nand NAND3 (N6407, N6404, N5786, N6028);
or OR2 (N6408, N6399, N1972);
not NOT1 (N6409, N6403);
buf BUF1 (N6410, N6406);
not NOT1 (N6411, N6374);
not NOT1 (N6412, N6380);
and AND3 (N6413, N6405, N5558, N3031);
nor NOR3 (N6414, N6408, N48, N3977);
nand NAND2 (N6415, N6414, N2287);
xor XOR2 (N6416, N6412, N6096);
endmodule