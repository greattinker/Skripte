// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13;

output N2983,N3008,N3006,N3003,N3011,N2996,N3012,N3010,N3005,N3013;

buf BUF1 (N14, N2);
nand NAND3 (N15, N8, N3, N10);
buf BUF1 (N16, N13);
and AND3 (N17, N3, N7, N3);
not NOT1 (N18, N16);
not NOT1 (N19, N9);
or OR2 (N20, N16, N4);
xor XOR2 (N21, N4, N15);
nand NAND2 (N22, N18, N20);
buf BUF1 (N23, N21);
and AND4 (N24, N19, N16, N23, N20);
nand NAND3 (N25, N5, N18, N11);
or OR3 (N26, N4, N5, N1);
not NOT1 (N27, N13);
nor NOR3 (N28, N23, N13, N19);
nand NAND4 (N29, N13, N23, N9, N3);
buf BUF1 (N30, N10);
and AND2 (N31, N14, N1);
nor NOR3 (N32, N17, N13, N12);
nand NAND4 (N33, N28, N11, N25, N19);
nor NOR2 (N34, N21, N24);
xor XOR2 (N35, N28, N2);
or OR4 (N36, N32, N2, N14, N20);
or OR3 (N37, N22, N12, N10);
xor XOR2 (N38, N35, N1);
buf BUF1 (N39, N30);
nand NAND2 (N40, N34, N11);
nor NOR4 (N41, N39, N22, N7, N39);
buf BUF1 (N42, N33);
or OR2 (N43, N41, N5);
nand NAND4 (N44, N43, N15, N1, N26);
not NOT1 (N45, N11);
buf BUF1 (N46, N29);
or OR2 (N47, N42, N9);
nor NOR3 (N48, N46, N8, N29);
buf BUF1 (N49, N27);
nand NAND2 (N50, N48, N3);
and AND2 (N51, N50, N35);
buf BUF1 (N52, N47);
and AND4 (N53, N45, N49, N26, N36);
or OR4 (N54, N13, N30, N23, N36);
and AND4 (N55, N25, N47, N54, N15);
or OR3 (N56, N13, N28, N45);
and AND2 (N57, N38, N54);
nand NAND3 (N58, N44, N41, N22);
nor NOR3 (N59, N52, N12, N39);
xor XOR2 (N60, N55, N6);
or OR4 (N61, N53, N48, N31, N59);
or OR3 (N62, N54, N29, N10);
nand NAND2 (N63, N58, N3);
or OR4 (N64, N26, N44, N54, N44);
not NOT1 (N65, N57);
or OR3 (N66, N61, N33, N31);
and AND3 (N67, N51, N15, N19);
and AND3 (N68, N40, N20, N10);
nand NAND2 (N69, N63, N20);
and AND3 (N70, N60, N58, N57);
nand NAND3 (N71, N68, N33, N32);
not NOT1 (N72, N67);
not NOT1 (N73, N65);
not NOT1 (N74, N72);
not NOT1 (N75, N73);
or OR4 (N76, N66, N10, N61, N4);
or OR2 (N77, N76, N73);
or OR2 (N78, N56, N5);
and AND2 (N79, N64, N44);
xor XOR2 (N80, N77, N24);
nor NOR4 (N81, N69, N56, N14, N45);
not NOT1 (N82, N74);
nor NOR4 (N83, N62, N19, N46, N55);
not NOT1 (N84, N71);
xor XOR2 (N85, N75, N23);
nand NAND3 (N86, N80, N79, N31);
nor NOR2 (N87, N9, N19);
not NOT1 (N88, N86);
not NOT1 (N89, N78);
not NOT1 (N90, N85);
and AND4 (N91, N88, N88, N15, N55);
not NOT1 (N92, N91);
xor XOR2 (N93, N90, N10);
and AND4 (N94, N93, N49, N30, N77);
or OR2 (N95, N92, N37);
nor NOR4 (N96, N90, N3, N70, N54);
nand NAND2 (N97, N39, N42);
and AND3 (N98, N95, N12, N46);
or OR2 (N99, N98, N88);
not NOT1 (N100, N99);
nor NOR4 (N101, N81, N50, N98, N68);
nor NOR4 (N102, N82, N98, N20, N84);
nand NAND2 (N103, N101, N53);
buf BUF1 (N104, N12);
and AND4 (N105, N83, N5, N65, N79);
nand NAND3 (N106, N97, N86, N29);
not NOT1 (N107, N103);
or OR3 (N108, N94, N87, N67);
xor XOR2 (N109, N102, N16);
nor NOR4 (N110, N16, N42, N92, N42);
xor XOR2 (N111, N89, N86);
or OR3 (N112, N107, N6, N79);
not NOT1 (N113, N108);
xor XOR2 (N114, N111, N74);
and AND4 (N115, N110, N37, N28, N68);
not NOT1 (N116, N106);
and AND3 (N117, N115, N104, N84);
or OR2 (N118, N63, N117);
buf BUF1 (N119, N98);
nor NOR3 (N120, N109, N57, N30);
or OR3 (N121, N113, N41, N42);
not NOT1 (N122, N118);
not NOT1 (N123, N121);
xor XOR2 (N124, N105, N90);
buf BUF1 (N125, N123);
not NOT1 (N126, N119);
not NOT1 (N127, N124);
or OR2 (N128, N114, N85);
nand NAND3 (N129, N120, N43, N33);
buf BUF1 (N130, N126);
xor XOR2 (N131, N100, N28);
and AND3 (N132, N116, N78, N2);
and AND2 (N133, N127, N131);
nand NAND3 (N134, N58, N70, N22);
and AND3 (N135, N132, N128, N71);
and AND2 (N136, N130, N133);
not NOT1 (N137, N14);
or OR3 (N138, N82, N134, N81);
not NOT1 (N139, N113);
buf BUF1 (N140, N136);
and AND4 (N141, N140, N107, N49, N18);
not NOT1 (N142, N137);
nand NAND2 (N143, N129, N87);
nor NOR4 (N144, N112, N111, N1, N72);
nor NOR2 (N145, N125, N76);
and AND4 (N146, N145, N98, N61, N133);
buf BUF1 (N147, N135);
nor NOR4 (N148, N146, N1, N71, N63);
and AND3 (N149, N139, N83, N67);
or OR4 (N150, N143, N4, N94, N26);
and AND3 (N151, N147, N16, N97);
nand NAND2 (N152, N144, N28);
not NOT1 (N153, N122);
xor XOR2 (N154, N150, N52);
nor NOR2 (N155, N149, N125);
and AND2 (N156, N138, N25);
nor NOR2 (N157, N155, N140);
xor XOR2 (N158, N152, N38);
buf BUF1 (N159, N96);
buf BUF1 (N160, N142);
not NOT1 (N161, N158);
not NOT1 (N162, N161);
and AND3 (N163, N162, N152, N52);
xor XOR2 (N164, N160, N59);
nor NOR3 (N165, N151, N15, N77);
nand NAND2 (N166, N164, N52);
buf BUF1 (N167, N163);
or OR3 (N168, N148, N6, N127);
or OR3 (N169, N165, N89, N112);
not NOT1 (N170, N156);
not NOT1 (N171, N169);
buf BUF1 (N172, N168);
buf BUF1 (N173, N157);
xor XOR2 (N174, N172, N131);
or OR3 (N175, N174, N43, N60);
not NOT1 (N176, N154);
and AND4 (N177, N159, N42, N175, N61);
and AND2 (N178, N117, N117);
xor XOR2 (N179, N141, N59);
xor XOR2 (N180, N176, N145);
xor XOR2 (N181, N179, N98);
and AND3 (N182, N153, N56, N15);
nand NAND4 (N183, N182, N97, N42, N133);
nand NAND2 (N184, N173, N163);
not NOT1 (N185, N166);
xor XOR2 (N186, N178, N67);
and AND4 (N187, N177, N162, N161, N179);
nor NOR3 (N188, N184, N51, N152);
xor XOR2 (N189, N171, N28);
buf BUF1 (N190, N170);
or OR4 (N191, N188, N125, N76, N181);
not NOT1 (N192, N73);
not NOT1 (N193, N189);
or OR2 (N194, N193, N74);
not NOT1 (N195, N192);
nor NOR4 (N196, N183, N144, N141, N78);
or OR3 (N197, N167, N126, N120);
nor NOR4 (N198, N196, N133, N163, N75);
nor NOR2 (N199, N198, N120);
nor NOR2 (N200, N195, N95);
and AND2 (N201, N185, N23);
xor XOR2 (N202, N194, N33);
and AND2 (N203, N199, N70);
xor XOR2 (N204, N202, N21);
xor XOR2 (N205, N187, N91);
not NOT1 (N206, N203);
xor XOR2 (N207, N197, N174);
or OR3 (N208, N180, N22, N78);
xor XOR2 (N209, N191, N145);
not NOT1 (N210, N204);
and AND4 (N211, N186, N129, N185, N140);
nand NAND3 (N212, N190, N186, N185);
xor XOR2 (N213, N206, N109);
nand NAND2 (N214, N211, N134);
and AND2 (N215, N210, N187);
buf BUF1 (N216, N205);
nor NOR4 (N217, N201, N26, N202, N209);
buf BUF1 (N218, N214);
or OR3 (N219, N30, N123, N183);
buf BUF1 (N220, N207);
xor XOR2 (N221, N212, N74);
or OR4 (N222, N220, N213, N214, N30);
buf BUF1 (N223, N192);
nand NAND2 (N224, N208, N10);
nor NOR4 (N225, N216, N224, N109, N171);
or OR3 (N226, N31, N201, N39);
not NOT1 (N227, N226);
xor XOR2 (N228, N217, N112);
nand NAND2 (N229, N225, N93);
xor XOR2 (N230, N228, N40);
or OR3 (N231, N230, N151, N128);
or OR2 (N232, N222, N52);
nand NAND4 (N233, N219, N20, N52, N133);
xor XOR2 (N234, N227, N188);
xor XOR2 (N235, N218, N217);
nor NOR4 (N236, N231, N178, N58, N223);
xor XOR2 (N237, N181, N24);
or OR2 (N238, N236, N140);
buf BUF1 (N239, N221);
buf BUF1 (N240, N237);
buf BUF1 (N241, N238);
nor NOR2 (N242, N240, N122);
xor XOR2 (N243, N233, N164);
xor XOR2 (N244, N234, N218);
nor NOR3 (N245, N232, N1, N231);
and AND2 (N246, N235, N22);
and AND3 (N247, N243, N240, N5);
buf BUF1 (N248, N200);
nand NAND3 (N249, N229, N197, N13);
nor NOR4 (N250, N245, N87, N196, N183);
and AND2 (N251, N247, N148);
and AND4 (N252, N241, N241, N127, N194);
nor NOR4 (N253, N215, N84, N144, N212);
or OR3 (N254, N244, N178, N52);
xor XOR2 (N255, N254, N148);
and AND2 (N256, N239, N222);
xor XOR2 (N257, N246, N21);
buf BUF1 (N258, N252);
buf BUF1 (N259, N251);
buf BUF1 (N260, N248);
nor NOR4 (N261, N260, N66, N118, N85);
nand NAND3 (N262, N258, N45, N2);
xor XOR2 (N263, N256, N53);
not NOT1 (N264, N249);
nor NOR4 (N265, N257, N181, N182, N191);
or OR2 (N266, N255, N23);
and AND4 (N267, N242, N230, N106, N174);
buf BUF1 (N268, N264);
and AND2 (N269, N250, N175);
buf BUF1 (N270, N265);
nand NAND4 (N271, N261, N77, N60, N100);
nor NOR3 (N272, N259, N199, N217);
or OR4 (N273, N253, N135, N148, N155);
and AND2 (N274, N268, N166);
and AND2 (N275, N262, N250);
nor NOR4 (N276, N267, N241, N12, N231);
xor XOR2 (N277, N269, N245);
nor NOR3 (N278, N271, N146, N102);
nand NAND4 (N279, N278, N57, N115, N132);
xor XOR2 (N280, N272, N59);
xor XOR2 (N281, N266, N23);
buf BUF1 (N282, N281);
and AND4 (N283, N270, N198, N47, N12);
or OR2 (N284, N280, N77);
and AND3 (N285, N277, N1, N190);
buf BUF1 (N286, N273);
or OR4 (N287, N284, N179, N277, N19);
xor XOR2 (N288, N276, N271);
or OR3 (N289, N263, N185, N140);
xor XOR2 (N290, N274, N89);
nand NAND3 (N291, N282, N143, N188);
buf BUF1 (N292, N291);
nand NAND3 (N293, N287, N191, N264);
xor XOR2 (N294, N283, N49);
or OR2 (N295, N293, N208);
xor XOR2 (N296, N286, N233);
not NOT1 (N297, N289);
nand NAND4 (N298, N297, N173, N19, N244);
and AND4 (N299, N275, N298, N233, N257);
buf BUF1 (N300, N143);
or OR4 (N301, N300, N6, N25, N124);
xor XOR2 (N302, N299, N61);
and AND3 (N303, N294, N223, N18);
and AND4 (N304, N302, N283, N201, N120);
nor NOR2 (N305, N304, N139);
nor NOR2 (N306, N303, N282);
nor NOR2 (N307, N301, N155);
nor NOR2 (N308, N290, N82);
buf BUF1 (N309, N307);
xor XOR2 (N310, N279, N156);
not NOT1 (N311, N296);
or OR2 (N312, N311, N205);
nand NAND4 (N313, N306, N309, N144, N144);
buf BUF1 (N314, N60);
nor NOR4 (N315, N314, N144, N179, N47);
not NOT1 (N316, N292);
and AND2 (N317, N316, N277);
xor XOR2 (N318, N317, N57);
xor XOR2 (N319, N315, N59);
nand NAND4 (N320, N288, N255, N120, N289);
buf BUF1 (N321, N320);
not NOT1 (N322, N321);
or OR4 (N323, N322, N287, N113, N56);
xor XOR2 (N324, N305, N230);
buf BUF1 (N325, N285);
not NOT1 (N326, N325);
not NOT1 (N327, N313);
not NOT1 (N328, N295);
nor NOR3 (N329, N326, N315, N53);
nand NAND4 (N330, N319, N6, N115, N179);
xor XOR2 (N331, N312, N128);
nand NAND2 (N332, N329, N244);
buf BUF1 (N333, N310);
and AND4 (N334, N324, N241, N149, N156);
buf BUF1 (N335, N333);
or OR2 (N336, N332, N51);
or OR2 (N337, N330, N249);
buf BUF1 (N338, N318);
not NOT1 (N339, N323);
not NOT1 (N340, N308);
and AND3 (N341, N335, N189, N49);
and AND4 (N342, N341, N250, N326, N171);
buf BUF1 (N343, N334);
not NOT1 (N344, N331);
buf BUF1 (N345, N344);
nand NAND3 (N346, N337, N286, N200);
and AND2 (N347, N342, N78);
not NOT1 (N348, N345);
and AND4 (N349, N348, N126, N139, N344);
not NOT1 (N350, N338);
not NOT1 (N351, N349);
or OR2 (N352, N340, N291);
nor NOR3 (N353, N343, N34, N137);
or OR2 (N354, N328, N139);
or OR2 (N355, N327, N248);
buf BUF1 (N356, N350);
nor NOR4 (N357, N347, N332, N281, N187);
or OR2 (N358, N352, N284);
nor NOR2 (N359, N356, N180);
buf BUF1 (N360, N336);
not NOT1 (N361, N354);
nand NAND2 (N362, N346, N361);
nand NAND3 (N363, N320, N322, N304);
nand NAND3 (N364, N363, N348, N355);
nor NOR4 (N365, N203, N331, N299, N12);
xor XOR2 (N366, N351, N272);
or OR4 (N367, N360, N192, N198, N210);
nand NAND3 (N368, N362, N212, N307);
and AND4 (N369, N353, N144, N24, N352);
xor XOR2 (N370, N369, N115);
or OR2 (N371, N359, N232);
or OR2 (N372, N357, N242);
not NOT1 (N373, N370);
buf BUF1 (N374, N339);
not NOT1 (N375, N365);
xor XOR2 (N376, N375, N338);
nand NAND2 (N377, N372, N290);
nor NOR3 (N378, N371, N167, N108);
nand NAND4 (N379, N377, N149, N320, N42);
not NOT1 (N380, N376);
or OR3 (N381, N373, N228, N186);
and AND3 (N382, N366, N167, N25);
and AND4 (N383, N374, N76, N307, N326);
xor XOR2 (N384, N358, N246);
or OR3 (N385, N379, N124, N268);
or OR4 (N386, N385, N105, N320, N69);
or OR2 (N387, N386, N168);
nand NAND4 (N388, N378, N266, N142, N90);
xor XOR2 (N389, N368, N40);
nand NAND2 (N390, N364, N32);
not NOT1 (N391, N367);
xor XOR2 (N392, N390, N23);
nand NAND4 (N393, N391, N42, N278, N378);
nor NOR4 (N394, N384, N182, N318, N238);
and AND2 (N395, N387, N279);
or OR2 (N396, N389, N355);
nor NOR3 (N397, N394, N221, N153);
xor XOR2 (N398, N392, N265);
nor NOR2 (N399, N383, N160);
or OR2 (N400, N399, N207);
or OR2 (N401, N397, N19);
buf BUF1 (N402, N380);
or OR3 (N403, N400, N277, N339);
nor NOR4 (N404, N393, N32, N242, N5);
buf BUF1 (N405, N396);
xor XOR2 (N406, N398, N325);
not NOT1 (N407, N388);
and AND3 (N408, N405, N279, N303);
nand NAND2 (N409, N404, N292);
or OR3 (N410, N407, N341, N191);
nand NAND3 (N411, N403, N32, N237);
nor NOR2 (N412, N402, N242);
xor XOR2 (N413, N408, N141);
buf BUF1 (N414, N395);
nand NAND3 (N415, N382, N230, N220);
or OR2 (N416, N406, N274);
buf BUF1 (N417, N413);
and AND2 (N418, N401, N126);
or OR4 (N419, N409, N195, N170, N125);
not NOT1 (N420, N381);
nand NAND3 (N421, N410, N78, N100);
nor NOR2 (N422, N411, N57);
nand NAND4 (N423, N415, N212, N39, N59);
or OR4 (N424, N422, N404, N133, N90);
not NOT1 (N425, N414);
xor XOR2 (N426, N425, N380);
nand NAND3 (N427, N424, N212, N243);
xor XOR2 (N428, N416, N198);
or OR2 (N429, N421, N428);
nand NAND2 (N430, N21, N25);
and AND3 (N431, N430, N10, N333);
xor XOR2 (N432, N429, N358);
or OR3 (N433, N417, N53, N84);
or OR2 (N434, N432, N173);
xor XOR2 (N435, N420, N283);
not NOT1 (N436, N423);
nand NAND4 (N437, N426, N235, N351, N36);
buf BUF1 (N438, N436);
or OR4 (N439, N434, N387, N166, N341);
or OR2 (N440, N433, N109);
nor NOR2 (N441, N437, N390);
xor XOR2 (N442, N435, N85);
and AND2 (N443, N419, N342);
not NOT1 (N444, N431);
not NOT1 (N445, N427);
xor XOR2 (N446, N441, N189);
nor NOR4 (N447, N412, N6, N50, N293);
not NOT1 (N448, N445);
buf BUF1 (N449, N443);
nand NAND4 (N450, N448, N277, N351, N2);
nor NOR4 (N451, N440, N66, N194, N110);
or OR3 (N452, N438, N360, N343);
nor NOR4 (N453, N446, N75, N325, N157);
and AND4 (N454, N447, N213, N293, N435);
nor NOR4 (N455, N454, N263, N123, N414);
nand NAND4 (N456, N449, N430, N134, N64);
or OR2 (N457, N455, N30);
xor XOR2 (N458, N457, N226);
nand NAND4 (N459, N450, N189, N199, N17);
buf BUF1 (N460, N444);
not NOT1 (N461, N418);
nor NOR2 (N462, N456, N8);
buf BUF1 (N463, N462);
nand NAND3 (N464, N459, N71, N153);
not NOT1 (N465, N442);
or OR3 (N466, N452, N182, N18);
xor XOR2 (N467, N461, N231);
nand NAND3 (N468, N463, N57, N394);
nor NOR3 (N469, N453, N293, N421);
buf BUF1 (N470, N460);
and AND3 (N471, N467, N306, N341);
not NOT1 (N472, N451);
nand NAND2 (N473, N471, N306);
nor NOR3 (N474, N465, N13, N26);
and AND4 (N475, N473, N175, N269, N263);
nand NAND2 (N476, N475, N364);
or OR3 (N477, N470, N102, N447);
nand NAND3 (N478, N477, N428, N133);
buf BUF1 (N479, N468);
nor NOR2 (N480, N464, N81);
and AND2 (N481, N474, N24);
xor XOR2 (N482, N472, N131);
nand NAND2 (N483, N482, N313);
nor NOR2 (N484, N481, N135);
buf BUF1 (N485, N483);
not NOT1 (N486, N466);
not NOT1 (N487, N478);
xor XOR2 (N488, N439, N189);
nor NOR3 (N489, N485, N346, N113);
not NOT1 (N490, N480);
buf BUF1 (N491, N469);
nand NAND3 (N492, N458, N348, N444);
and AND3 (N493, N489, N485, N83);
nand NAND4 (N494, N476, N155, N254, N259);
xor XOR2 (N495, N479, N109);
not NOT1 (N496, N488);
nor NOR2 (N497, N495, N258);
buf BUF1 (N498, N484);
and AND2 (N499, N497, N466);
or OR4 (N500, N492, N290, N325, N167);
buf BUF1 (N501, N496);
nand NAND2 (N502, N500, N155);
buf BUF1 (N503, N499);
nor NOR3 (N504, N486, N112, N241);
xor XOR2 (N505, N493, N399);
xor XOR2 (N506, N494, N50);
buf BUF1 (N507, N506);
nor NOR2 (N508, N505, N429);
xor XOR2 (N509, N508, N77);
or OR4 (N510, N509, N171, N311, N217);
buf BUF1 (N511, N501);
buf BUF1 (N512, N498);
and AND2 (N513, N512, N369);
nand NAND4 (N514, N510, N149, N211, N472);
not NOT1 (N515, N503);
and AND3 (N516, N514, N444, N483);
nor NOR2 (N517, N511, N77);
nand NAND4 (N518, N507, N330, N65, N12);
xor XOR2 (N519, N487, N323);
nor NOR2 (N520, N516, N467);
xor XOR2 (N521, N518, N164);
xor XOR2 (N522, N491, N484);
nand NAND4 (N523, N521, N150, N138, N481);
xor XOR2 (N524, N513, N84);
not NOT1 (N525, N490);
nand NAND3 (N526, N525, N31, N105);
xor XOR2 (N527, N523, N354);
or OR3 (N528, N522, N284, N330);
or OR4 (N529, N517, N357, N485, N43);
and AND2 (N530, N524, N428);
nand NAND4 (N531, N515, N365, N171, N340);
nand NAND3 (N532, N504, N59, N94);
not NOT1 (N533, N528);
and AND4 (N534, N532, N509, N470, N358);
nor NOR2 (N535, N520, N230);
and AND3 (N536, N526, N35, N494);
nand NAND4 (N537, N531, N425, N531, N130);
xor XOR2 (N538, N536, N501);
nand NAND2 (N539, N533, N88);
xor XOR2 (N540, N539, N242);
not NOT1 (N541, N537);
not NOT1 (N542, N535);
not NOT1 (N543, N534);
nand NAND3 (N544, N543, N534, N391);
xor XOR2 (N545, N529, N110);
and AND4 (N546, N544, N421, N164, N312);
or OR3 (N547, N527, N334, N406);
nor NOR3 (N548, N502, N486, N409);
and AND4 (N549, N545, N411, N120, N468);
nor NOR4 (N550, N542, N385, N27, N442);
nand NAND4 (N551, N538, N380, N390, N275);
buf BUF1 (N552, N547);
buf BUF1 (N553, N548);
nand NAND2 (N554, N550, N511);
nor NOR2 (N555, N541, N43);
nor NOR3 (N556, N530, N401, N383);
xor XOR2 (N557, N555, N459);
nand NAND3 (N558, N557, N305, N168);
or OR4 (N559, N540, N380, N547, N457);
or OR2 (N560, N558, N117);
or OR4 (N561, N556, N325, N181, N130);
and AND2 (N562, N519, N254);
and AND3 (N563, N562, N478, N449);
nor NOR4 (N564, N549, N482, N85, N62);
xor XOR2 (N565, N561, N268);
nand NAND3 (N566, N563, N208, N446);
buf BUF1 (N567, N551);
buf BUF1 (N568, N553);
not NOT1 (N569, N567);
nor NOR4 (N570, N565, N410, N51, N510);
not NOT1 (N571, N546);
and AND4 (N572, N560, N43, N287, N127);
nand NAND2 (N573, N564, N355);
buf BUF1 (N574, N568);
not NOT1 (N575, N566);
not NOT1 (N576, N569);
or OR2 (N577, N554, N29);
buf BUF1 (N578, N552);
buf BUF1 (N579, N576);
not NOT1 (N580, N574);
or OR3 (N581, N559, N57, N180);
and AND4 (N582, N573, N208, N275, N31);
or OR2 (N583, N571, N432);
xor XOR2 (N584, N575, N503);
buf BUF1 (N585, N570);
xor XOR2 (N586, N578, N469);
nand NAND2 (N587, N583, N388);
buf BUF1 (N588, N582);
or OR4 (N589, N579, N99, N358, N82);
nor NOR4 (N590, N577, N55, N220, N507);
buf BUF1 (N591, N587);
xor XOR2 (N592, N581, N119);
nor NOR2 (N593, N589, N452);
and AND3 (N594, N572, N31, N51);
buf BUF1 (N595, N590);
xor XOR2 (N596, N592, N367);
nor NOR3 (N597, N591, N107, N271);
buf BUF1 (N598, N593);
nor NOR4 (N599, N598, N16, N475, N284);
or OR3 (N600, N597, N141, N456);
not NOT1 (N601, N594);
nor NOR3 (N602, N584, N369, N578);
or OR3 (N603, N596, N298, N95);
xor XOR2 (N604, N586, N51);
nor NOR4 (N605, N588, N287, N217, N186);
not NOT1 (N606, N585);
not NOT1 (N607, N601);
nor NOR2 (N608, N606, N233);
buf BUF1 (N609, N605);
not NOT1 (N610, N580);
not NOT1 (N611, N608);
nand NAND4 (N612, N602, N302, N566, N472);
buf BUF1 (N613, N612);
xor XOR2 (N614, N599, N489);
buf BUF1 (N615, N611);
nand NAND3 (N616, N615, N222, N363);
nand NAND4 (N617, N610, N510, N335, N351);
buf BUF1 (N618, N617);
not NOT1 (N619, N613);
xor XOR2 (N620, N603, N107);
or OR2 (N621, N604, N555);
nand NAND2 (N622, N621, N558);
nor NOR2 (N623, N620, N147);
xor XOR2 (N624, N623, N118);
buf BUF1 (N625, N618);
nand NAND2 (N626, N622, N580);
and AND2 (N627, N624, N12);
and AND3 (N628, N600, N92, N257);
nor NOR2 (N629, N625, N331);
buf BUF1 (N630, N628);
nand NAND3 (N631, N629, N447, N107);
or OR3 (N632, N631, N608, N175);
buf BUF1 (N633, N595);
buf BUF1 (N634, N616);
xor XOR2 (N635, N619, N478);
and AND2 (N636, N634, N34);
or OR4 (N637, N636, N39, N9, N407);
xor XOR2 (N638, N635, N579);
or OR4 (N639, N633, N51, N338, N576);
or OR3 (N640, N626, N175, N85);
nand NAND2 (N641, N609, N638);
nor NOR4 (N642, N385, N568, N361, N638);
buf BUF1 (N643, N642);
nor NOR2 (N644, N614, N352);
not NOT1 (N645, N627);
buf BUF1 (N646, N607);
or OR2 (N647, N630, N517);
nand NAND3 (N648, N644, N490, N316);
xor XOR2 (N649, N646, N119);
or OR2 (N650, N639, N501);
or OR2 (N651, N650, N375);
and AND4 (N652, N643, N220, N63, N183);
and AND2 (N653, N651, N536);
xor XOR2 (N654, N645, N108);
or OR2 (N655, N641, N110);
xor XOR2 (N656, N652, N431);
not NOT1 (N657, N654);
xor XOR2 (N658, N648, N76);
and AND3 (N659, N632, N11, N64);
xor XOR2 (N660, N640, N139);
nor NOR3 (N661, N658, N231, N516);
nand NAND3 (N662, N649, N181, N192);
nand NAND3 (N663, N637, N357, N186);
xor XOR2 (N664, N647, N311);
not NOT1 (N665, N661);
nand NAND2 (N666, N662, N538);
and AND3 (N667, N659, N250, N619);
not NOT1 (N668, N653);
nor NOR4 (N669, N656, N5, N94, N394);
not NOT1 (N670, N665);
or OR4 (N671, N667, N385, N520, N433);
nor NOR2 (N672, N670, N24);
or OR2 (N673, N671, N368);
xor XOR2 (N674, N660, N356);
nor NOR4 (N675, N669, N254, N188, N280);
buf BUF1 (N676, N675);
nor NOR3 (N677, N674, N442, N238);
buf BUF1 (N678, N657);
not NOT1 (N679, N664);
nor NOR4 (N680, N678, N75, N547, N281);
nand NAND3 (N681, N666, N391, N75);
nor NOR3 (N682, N668, N190, N461);
not NOT1 (N683, N673);
or OR3 (N684, N676, N175, N131);
and AND2 (N685, N679, N112);
xor XOR2 (N686, N672, N499);
xor XOR2 (N687, N683, N5);
or OR4 (N688, N686, N304, N580, N342);
nand NAND4 (N689, N682, N651, N667, N431);
and AND2 (N690, N663, N576);
not NOT1 (N691, N687);
buf BUF1 (N692, N690);
or OR2 (N693, N655, N244);
not NOT1 (N694, N691);
nor NOR3 (N695, N680, N325, N96);
xor XOR2 (N696, N681, N89);
and AND3 (N697, N688, N305, N447);
nand NAND2 (N698, N684, N222);
not NOT1 (N699, N685);
nor NOR4 (N700, N696, N83, N431, N426);
not NOT1 (N701, N700);
nand NAND2 (N702, N692, N547);
buf BUF1 (N703, N693);
not NOT1 (N704, N701);
nand NAND2 (N705, N703, N506);
xor XOR2 (N706, N704, N455);
nor NOR4 (N707, N697, N115, N296, N484);
xor XOR2 (N708, N694, N375);
or OR4 (N709, N705, N73, N78, N628);
nor NOR2 (N710, N689, N452);
buf BUF1 (N711, N677);
nand NAND3 (N712, N709, N336, N72);
and AND4 (N713, N708, N667, N251, N501);
or OR3 (N714, N702, N206, N238);
not NOT1 (N715, N695);
buf BUF1 (N716, N706);
nand NAND4 (N717, N715, N600, N109, N577);
nand NAND2 (N718, N716, N329);
xor XOR2 (N719, N710, N28);
buf BUF1 (N720, N718);
nor NOR2 (N721, N717, N99);
not NOT1 (N722, N699);
xor XOR2 (N723, N719, N646);
nand NAND3 (N724, N712, N166, N279);
nand NAND4 (N725, N721, N574, N263, N461);
xor XOR2 (N726, N723, N681);
and AND2 (N727, N698, N634);
nor NOR4 (N728, N724, N486, N709, N393);
not NOT1 (N729, N714);
buf BUF1 (N730, N728);
not NOT1 (N731, N722);
nor NOR4 (N732, N707, N583, N573, N728);
nand NAND4 (N733, N729, N486, N58, N429);
or OR4 (N734, N726, N469, N598, N349);
nor NOR4 (N735, N720, N306, N600, N399);
not NOT1 (N736, N713);
xor XOR2 (N737, N732, N170);
not NOT1 (N738, N737);
xor XOR2 (N739, N734, N719);
not NOT1 (N740, N730);
xor XOR2 (N741, N725, N416);
buf BUF1 (N742, N736);
and AND4 (N743, N738, N186, N664, N342);
not NOT1 (N744, N733);
or OR3 (N745, N731, N124, N697);
nand NAND2 (N746, N744, N385);
buf BUF1 (N747, N742);
nand NAND2 (N748, N735, N482);
not NOT1 (N749, N743);
not NOT1 (N750, N741);
not NOT1 (N751, N750);
or OR3 (N752, N727, N177, N367);
xor XOR2 (N753, N739, N701);
xor XOR2 (N754, N751, N138);
or OR4 (N755, N754, N271, N526, N166);
xor XOR2 (N756, N753, N535);
and AND4 (N757, N747, N72, N403, N129);
nand NAND3 (N758, N746, N668, N66);
nand NAND3 (N759, N758, N194, N229);
nor NOR3 (N760, N740, N205, N578);
nand NAND2 (N761, N749, N649);
or OR3 (N762, N756, N63, N484);
nor NOR3 (N763, N759, N233, N43);
not NOT1 (N764, N761);
buf BUF1 (N765, N760);
nor NOR4 (N766, N711, N613, N141, N717);
nor NOR3 (N767, N748, N141, N183);
buf BUF1 (N768, N764);
not NOT1 (N769, N762);
nor NOR3 (N770, N745, N493, N405);
buf BUF1 (N771, N755);
buf BUF1 (N772, N769);
nor NOR4 (N773, N763, N502, N280, N44);
buf BUF1 (N774, N767);
nand NAND3 (N775, N770, N413, N580);
xor XOR2 (N776, N774, N724);
and AND2 (N777, N776, N88);
and AND3 (N778, N771, N184, N61);
or OR4 (N779, N768, N246, N577, N552);
and AND3 (N780, N778, N260, N176);
nand NAND4 (N781, N777, N186, N340, N196);
and AND2 (N782, N781, N471);
buf BUF1 (N783, N775);
xor XOR2 (N784, N782, N623);
and AND4 (N785, N784, N629, N619, N245);
nand NAND4 (N786, N785, N393, N547, N593);
not NOT1 (N787, N773);
or OR3 (N788, N752, N519, N768);
buf BUF1 (N789, N779);
nor NOR3 (N790, N772, N454, N298);
and AND2 (N791, N780, N499);
not NOT1 (N792, N765);
nand NAND2 (N793, N792, N638);
xor XOR2 (N794, N787, N150);
or OR3 (N795, N793, N772, N661);
and AND3 (N796, N791, N67, N762);
and AND3 (N797, N796, N125, N383);
nor NOR3 (N798, N790, N630, N693);
and AND3 (N799, N783, N451, N80);
not NOT1 (N800, N798);
xor XOR2 (N801, N757, N554);
and AND2 (N802, N766, N117);
not NOT1 (N803, N788);
buf BUF1 (N804, N795);
and AND4 (N805, N789, N798, N566, N354);
and AND3 (N806, N786, N214, N409);
not NOT1 (N807, N802);
nor NOR2 (N808, N794, N155);
nor NOR3 (N809, N803, N421, N413);
not NOT1 (N810, N801);
or OR4 (N811, N809, N406, N571, N565);
or OR3 (N812, N800, N18, N213);
buf BUF1 (N813, N811);
and AND3 (N814, N813, N609, N460);
xor XOR2 (N815, N805, N381);
xor XOR2 (N816, N806, N637);
or OR2 (N817, N804, N462);
and AND4 (N818, N817, N231, N156, N521);
xor XOR2 (N819, N797, N323);
not NOT1 (N820, N814);
not NOT1 (N821, N808);
and AND4 (N822, N812, N398, N640, N7);
nor NOR2 (N823, N818, N111);
or OR2 (N824, N821, N567);
and AND3 (N825, N822, N726, N634);
buf BUF1 (N826, N816);
not NOT1 (N827, N823);
nor NOR3 (N828, N826, N210, N605);
not NOT1 (N829, N824);
xor XOR2 (N830, N827, N236);
not NOT1 (N831, N830);
buf BUF1 (N832, N799);
or OR2 (N833, N828, N549);
or OR2 (N834, N832, N113);
nor NOR4 (N835, N833, N512, N781, N665);
or OR2 (N836, N835, N791);
buf BUF1 (N837, N815);
or OR3 (N838, N829, N748, N116);
nor NOR3 (N839, N831, N379, N91);
buf BUF1 (N840, N838);
nand NAND4 (N841, N834, N440, N145, N92);
not NOT1 (N842, N839);
xor XOR2 (N843, N819, N658);
nor NOR3 (N844, N837, N176, N745);
nor NOR4 (N845, N844, N449, N549, N197);
or OR3 (N846, N820, N206, N695);
and AND4 (N847, N810, N386, N142, N117);
nor NOR3 (N848, N825, N171, N187);
and AND3 (N849, N840, N520, N811);
buf BUF1 (N850, N843);
and AND4 (N851, N836, N818, N373, N635);
nor NOR3 (N852, N841, N804, N767);
not NOT1 (N853, N845);
not NOT1 (N854, N847);
and AND3 (N855, N852, N285, N103);
or OR4 (N856, N807, N290, N626, N343);
not NOT1 (N857, N856);
nor NOR4 (N858, N857, N118, N621, N283);
or OR2 (N859, N850, N345);
xor XOR2 (N860, N848, N811);
or OR4 (N861, N846, N397, N753, N463);
buf BUF1 (N862, N854);
buf BUF1 (N863, N861);
or OR4 (N864, N851, N516, N249, N51);
or OR3 (N865, N862, N323, N847);
or OR3 (N866, N855, N178, N617);
nor NOR4 (N867, N859, N823, N691, N8);
and AND2 (N868, N842, N725);
nand NAND3 (N869, N863, N353, N672);
or OR4 (N870, N868, N139, N122, N677);
or OR4 (N871, N865, N507, N343, N304);
xor XOR2 (N872, N867, N613);
and AND2 (N873, N869, N423);
nor NOR3 (N874, N864, N138, N78);
nand NAND2 (N875, N873, N124);
or OR3 (N876, N866, N864, N752);
not NOT1 (N877, N871);
nand NAND3 (N878, N858, N556, N789);
xor XOR2 (N879, N874, N97);
not NOT1 (N880, N853);
or OR4 (N881, N877, N288, N92, N764);
buf BUF1 (N882, N879);
nor NOR2 (N883, N870, N690);
not NOT1 (N884, N881);
not NOT1 (N885, N876);
not NOT1 (N886, N880);
nor NOR4 (N887, N872, N141, N270, N111);
not NOT1 (N888, N887);
not NOT1 (N889, N860);
not NOT1 (N890, N849);
buf BUF1 (N891, N878);
not NOT1 (N892, N882);
nand NAND3 (N893, N889, N835, N594);
buf BUF1 (N894, N884);
buf BUF1 (N895, N894);
nand NAND4 (N896, N892, N807, N573, N260);
buf BUF1 (N897, N888);
buf BUF1 (N898, N893);
and AND4 (N899, N898, N360, N342, N868);
nand NAND2 (N900, N896, N788);
and AND4 (N901, N897, N736, N668, N701);
or OR3 (N902, N891, N247, N502);
buf BUF1 (N903, N875);
and AND2 (N904, N895, N182);
or OR2 (N905, N885, N289);
or OR4 (N906, N904, N250, N855, N715);
nor NOR4 (N907, N901, N133, N369, N825);
or OR2 (N908, N890, N675);
xor XOR2 (N909, N907, N403);
nor NOR3 (N910, N900, N870, N572);
buf BUF1 (N911, N883);
nand NAND2 (N912, N902, N462);
xor XOR2 (N913, N908, N283);
xor XOR2 (N914, N905, N94);
xor XOR2 (N915, N906, N138);
and AND3 (N916, N903, N719, N436);
and AND2 (N917, N910, N784);
nand NAND4 (N918, N917, N799, N823, N249);
or OR3 (N919, N914, N535, N335);
buf BUF1 (N920, N899);
or OR2 (N921, N909, N376);
and AND4 (N922, N886, N813, N570, N16);
not NOT1 (N923, N913);
not NOT1 (N924, N922);
buf BUF1 (N925, N921);
xor XOR2 (N926, N923, N643);
or OR4 (N927, N924, N844, N824, N40);
or OR4 (N928, N915, N546, N365, N759);
nor NOR3 (N929, N925, N606, N413);
buf BUF1 (N930, N929);
xor XOR2 (N931, N927, N676);
or OR4 (N932, N919, N872, N385, N505);
not NOT1 (N933, N930);
and AND4 (N934, N928, N576, N667, N453);
or OR4 (N935, N912, N467, N722, N45);
nand NAND3 (N936, N911, N314, N393);
buf BUF1 (N937, N926);
or OR2 (N938, N918, N38);
xor XOR2 (N939, N935, N284);
and AND4 (N940, N938, N909, N268, N168);
nand NAND4 (N941, N939, N434, N564, N267);
nand NAND2 (N942, N941, N232);
not NOT1 (N943, N932);
xor XOR2 (N944, N933, N750);
nand NAND3 (N945, N931, N793, N456);
nand NAND2 (N946, N944, N583);
or OR3 (N947, N920, N802, N81);
or OR4 (N948, N946, N91, N767, N937);
not NOT1 (N949, N385);
and AND3 (N950, N949, N168, N862);
not NOT1 (N951, N950);
nor NOR3 (N952, N947, N65, N115);
nand NAND4 (N953, N943, N22, N91, N511);
or OR3 (N954, N916, N205, N322);
buf BUF1 (N955, N942);
xor XOR2 (N956, N945, N698);
xor XOR2 (N957, N955, N906);
and AND3 (N958, N940, N388, N805);
buf BUF1 (N959, N957);
or OR4 (N960, N958, N306, N267, N654);
nor NOR2 (N961, N953, N189);
xor XOR2 (N962, N934, N363);
or OR3 (N963, N962, N400, N474);
nor NOR2 (N964, N959, N559);
or OR3 (N965, N961, N446, N619);
xor XOR2 (N966, N956, N379);
or OR3 (N967, N965, N248, N911);
nand NAND4 (N968, N966, N413, N446, N384);
buf BUF1 (N969, N954);
and AND2 (N970, N963, N683);
nand NAND2 (N971, N936, N576);
nand NAND4 (N972, N951, N746, N665, N854);
nor NOR2 (N973, N964, N763);
and AND3 (N974, N973, N599, N879);
and AND4 (N975, N960, N802, N124, N18);
xor XOR2 (N976, N975, N360);
nand NAND2 (N977, N976, N568);
xor XOR2 (N978, N970, N219);
xor XOR2 (N979, N968, N537);
and AND4 (N980, N971, N446, N351, N192);
or OR3 (N981, N948, N594, N400);
and AND2 (N982, N978, N216);
or OR2 (N983, N972, N126);
nand NAND4 (N984, N983, N784, N176, N200);
nand NAND2 (N985, N967, N124);
nor NOR4 (N986, N979, N932, N130, N479);
nand NAND4 (N987, N977, N94, N61, N846);
or OR2 (N988, N987, N405);
nor NOR4 (N989, N969, N745, N616, N233);
nand NAND2 (N990, N952, N897);
and AND4 (N991, N989, N22, N553, N467);
not NOT1 (N992, N986);
nand NAND4 (N993, N988, N75, N135, N971);
nand NAND4 (N994, N984, N347, N498, N960);
nor NOR2 (N995, N981, N598);
nand NAND3 (N996, N982, N33, N505);
and AND3 (N997, N992, N396, N54);
nor NOR3 (N998, N995, N511, N929);
xor XOR2 (N999, N997, N813);
buf BUF1 (N1000, N974);
nor NOR4 (N1001, N998, N612, N378, N906);
not NOT1 (N1002, N980);
nand NAND3 (N1003, N993, N784, N183);
xor XOR2 (N1004, N991, N210);
or OR3 (N1005, N1001, N468, N742);
buf BUF1 (N1006, N999);
buf BUF1 (N1007, N1002);
xor XOR2 (N1008, N1007, N198);
xor XOR2 (N1009, N1006, N1008);
xor XOR2 (N1010, N462, N522);
nand NAND2 (N1011, N1010, N778);
xor XOR2 (N1012, N1005, N662);
nand NAND2 (N1013, N996, N289);
or OR2 (N1014, N1000, N126);
xor XOR2 (N1015, N994, N650);
and AND2 (N1016, N1003, N514);
and AND2 (N1017, N1015, N20);
and AND4 (N1018, N1016, N62, N416, N11);
or OR2 (N1019, N1009, N294);
nand NAND2 (N1020, N1017, N724);
not NOT1 (N1021, N1004);
or OR3 (N1022, N1021, N265, N792);
not NOT1 (N1023, N1019);
nand NAND4 (N1024, N1014, N624, N525, N138);
buf BUF1 (N1025, N1023);
buf BUF1 (N1026, N1025);
xor XOR2 (N1027, N985, N395);
nor NOR3 (N1028, N1022, N462, N105);
xor XOR2 (N1029, N1011, N483);
nand NAND3 (N1030, N1024, N458, N42);
nand NAND2 (N1031, N1029, N840);
or OR2 (N1032, N1031, N258);
buf BUF1 (N1033, N1032);
not NOT1 (N1034, N1033);
or OR3 (N1035, N1020, N937, N155);
and AND2 (N1036, N1028, N19);
or OR2 (N1037, N1026, N948);
nand NAND3 (N1038, N1012, N327, N890);
nor NOR3 (N1039, N1030, N345, N271);
buf BUF1 (N1040, N1018);
nand NAND2 (N1041, N1038, N712);
not NOT1 (N1042, N1013);
and AND3 (N1043, N990, N476, N297);
buf BUF1 (N1044, N1035);
not NOT1 (N1045, N1027);
not NOT1 (N1046, N1043);
and AND3 (N1047, N1037, N703, N499);
or OR4 (N1048, N1040, N321, N253, N437);
or OR3 (N1049, N1039, N701, N177);
and AND2 (N1050, N1045, N876);
not NOT1 (N1051, N1047);
xor XOR2 (N1052, N1042, N438);
nand NAND3 (N1053, N1049, N396, N705);
or OR2 (N1054, N1041, N641);
nor NOR4 (N1055, N1050, N54, N451, N331);
and AND3 (N1056, N1034, N999, N456);
or OR2 (N1057, N1056, N942);
not NOT1 (N1058, N1054);
not NOT1 (N1059, N1046);
and AND3 (N1060, N1036, N264, N585);
buf BUF1 (N1061, N1044);
not NOT1 (N1062, N1048);
buf BUF1 (N1063, N1051);
and AND2 (N1064, N1057, N165);
buf BUF1 (N1065, N1061);
buf BUF1 (N1066, N1065);
xor XOR2 (N1067, N1055, N362);
not NOT1 (N1068, N1058);
nand NAND3 (N1069, N1052, N1052, N662);
not NOT1 (N1070, N1062);
not NOT1 (N1071, N1067);
not NOT1 (N1072, N1071);
or OR4 (N1073, N1064, N641, N1045, N871);
buf BUF1 (N1074, N1069);
nor NOR3 (N1075, N1072, N654, N788);
or OR3 (N1076, N1068, N723, N816);
nand NAND2 (N1077, N1076, N547);
nor NOR3 (N1078, N1060, N324, N101);
buf BUF1 (N1079, N1075);
not NOT1 (N1080, N1063);
and AND3 (N1081, N1070, N445, N107);
nand NAND2 (N1082, N1081, N650);
or OR4 (N1083, N1080, N823, N388, N491);
xor XOR2 (N1084, N1066, N239);
not NOT1 (N1085, N1083);
not NOT1 (N1086, N1079);
nand NAND3 (N1087, N1053, N509, N268);
nand NAND3 (N1088, N1077, N1070, N841);
nor NOR3 (N1089, N1074, N822, N477);
and AND3 (N1090, N1089, N498, N842);
and AND3 (N1091, N1087, N548, N842);
or OR4 (N1092, N1073, N319, N746, N681);
buf BUF1 (N1093, N1090);
not NOT1 (N1094, N1084);
not NOT1 (N1095, N1088);
buf BUF1 (N1096, N1078);
buf BUF1 (N1097, N1093);
or OR3 (N1098, N1092, N49, N555);
or OR4 (N1099, N1094, N732, N610, N689);
nand NAND2 (N1100, N1099, N824);
and AND2 (N1101, N1100, N1029);
nor NOR3 (N1102, N1095, N593, N978);
nand NAND2 (N1103, N1101, N214);
xor XOR2 (N1104, N1091, N277);
buf BUF1 (N1105, N1082);
and AND3 (N1106, N1102, N783, N190);
nor NOR2 (N1107, N1106, N1015);
or OR4 (N1108, N1107, N303, N725, N113);
nor NOR3 (N1109, N1108, N234, N435);
xor XOR2 (N1110, N1105, N705);
xor XOR2 (N1111, N1085, N773);
or OR4 (N1112, N1104, N860, N385, N287);
and AND3 (N1113, N1112, N647, N56);
nor NOR3 (N1114, N1109, N194, N629);
or OR3 (N1115, N1103, N470, N453);
buf BUF1 (N1116, N1110);
xor XOR2 (N1117, N1113, N1007);
nand NAND2 (N1118, N1117, N1064);
not NOT1 (N1119, N1098);
not NOT1 (N1120, N1116);
nand NAND2 (N1121, N1120, N245);
and AND3 (N1122, N1115, N1034, N1064);
and AND3 (N1123, N1122, N921, N453);
not NOT1 (N1124, N1086);
nand NAND3 (N1125, N1059, N945, N52);
nand NAND2 (N1126, N1114, N670);
and AND3 (N1127, N1123, N680, N127);
not NOT1 (N1128, N1121);
and AND2 (N1129, N1126, N1118);
not NOT1 (N1130, N798);
not NOT1 (N1131, N1124);
nand NAND4 (N1132, N1111, N341, N782, N281);
xor XOR2 (N1133, N1125, N65);
xor XOR2 (N1134, N1127, N631);
xor XOR2 (N1135, N1096, N628);
nor NOR2 (N1136, N1132, N576);
or OR4 (N1137, N1136, N99, N872, N734);
nand NAND2 (N1138, N1135, N735);
buf BUF1 (N1139, N1119);
nand NAND3 (N1140, N1130, N493, N987);
not NOT1 (N1141, N1140);
or OR3 (N1142, N1128, N480, N486);
xor XOR2 (N1143, N1142, N793);
nor NOR4 (N1144, N1133, N253, N934, N371);
nor NOR3 (N1145, N1139, N101, N399);
and AND3 (N1146, N1138, N471, N670);
nor NOR3 (N1147, N1131, N358, N1060);
xor XOR2 (N1148, N1146, N1009);
xor XOR2 (N1149, N1145, N895);
xor XOR2 (N1150, N1141, N13);
nand NAND3 (N1151, N1149, N821, N861);
or OR2 (N1152, N1151, N541);
or OR4 (N1153, N1152, N1017, N289, N120);
buf BUF1 (N1154, N1134);
nor NOR3 (N1155, N1144, N419, N1135);
and AND4 (N1156, N1155, N577, N1110, N799);
and AND4 (N1157, N1156, N461, N696, N228);
not NOT1 (N1158, N1157);
buf BUF1 (N1159, N1129);
xor XOR2 (N1160, N1147, N585);
or OR3 (N1161, N1150, N15, N648);
nor NOR3 (N1162, N1097, N687, N950);
nor NOR4 (N1163, N1161, N595, N154, N108);
or OR3 (N1164, N1153, N68, N649);
not NOT1 (N1165, N1164);
nand NAND2 (N1166, N1154, N1153);
or OR3 (N1167, N1143, N44, N65);
xor XOR2 (N1168, N1165, N627);
nor NOR2 (N1169, N1148, N921);
nand NAND3 (N1170, N1166, N136, N707);
and AND3 (N1171, N1162, N20, N28);
and AND2 (N1172, N1160, N870);
xor XOR2 (N1173, N1159, N1047);
buf BUF1 (N1174, N1171);
or OR4 (N1175, N1137, N947, N551, N583);
nor NOR2 (N1176, N1158, N545);
buf BUF1 (N1177, N1167);
or OR2 (N1178, N1176, N520);
buf BUF1 (N1179, N1173);
nor NOR3 (N1180, N1169, N504, N900);
and AND3 (N1181, N1180, N143, N917);
not NOT1 (N1182, N1178);
nand NAND3 (N1183, N1182, N1, N200);
nor NOR4 (N1184, N1179, N699, N733, N871);
buf BUF1 (N1185, N1172);
and AND4 (N1186, N1185, N993, N940, N729);
or OR4 (N1187, N1184, N1094, N222, N177);
buf BUF1 (N1188, N1168);
nand NAND4 (N1189, N1163, N439, N379, N430);
and AND2 (N1190, N1189, N109);
buf BUF1 (N1191, N1188);
or OR4 (N1192, N1187, N139, N709, N1009);
and AND2 (N1193, N1181, N269);
and AND2 (N1194, N1177, N612);
or OR4 (N1195, N1170, N32, N66, N64);
nor NOR2 (N1196, N1174, N103);
nand NAND3 (N1197, N1195, N800, N36);
xor XOR2 (N1198, N1175, N886);
xor XOR2 (N1199, N1196, N619);
xor XOR2 (N1200, N1183, N479);
buf BUF1 (N1201, N1190);
not NOT1 (N1202, N1193);
or OR4 (N1203, N1201, N1033, N1007, N156);
and AND3 (N1204, N1191, N241, N440);
buf BUF1 (N1205, N1194);
xor XOR2 (N1206, N1203, N358);
xor XOR2 (N1207, N1192, N438);
not NOT1 (N1208, N1202);
xor XOR2 (N1209, N1204, N364);
buf BUF1 (N1210, N1209);
not NOT1 (N1211, N1200);
nor NOR3 (N1212, N1186, N920, N40);
or OR3 (N1213, N1199, N97, N1037);
not NOT1 (N1214, N1207);
nand NAND2 (N1215, N1208, N475);
or OR4 (N1216, N1197, N995, N392, N417);
and AND4 (N1217, N1212, N748, N764, N572);
not NOT1 (N1218, N1216);
nor NOR4 (N1219, N1217, N805, N586, N756);
and AND4 (N1220, N1205, N159, N428, N18);
nand NAND4 (N1221, N1211, N911, N489, N787);
not NOT1 (N1222, N1206);
nand NAND4 (N1223, N1214, N115, N1054, N781);
buf BUF1 (N1224, N1222);
nor NOR3 (N1225, N1221, N214, N130);
xor XOR2 (N1226, N1223, N1195);
not NOT1 (N1227, N1198);
nor NOR4 (N1228, N1227, N718, N848, N249);
nor NOR3 (N1229, N1210, N257, N31);
and AND2 (N1230, N1219, N1100);
nor NOR4 (N1231, N1229, N832, N1009, N336);
nand NAND2 (N1232, N1213, N444);
xor XOR2 (N1233, N1215, N137);
xor XOR2 (N1234, N1233, N767);
nand NAND2 (N1235, N1225, N1012);
xor XOR2 (N1236, N1224, N1166);
nand NAND4 (N1237, N1235, N782, N71, N463);
nor NOR3 (N1238, N1220, N835, N127);
not NOT1 (N1239, N1238);
or OR2 (N1240, N1230, N908);
and AND4 (N1241, N1232, N670, N960, N1200);
or OR2 (N1242, N1231, N240);
xor XOR2 (N1243, N1241, N51);
xor XOR2 (N1244, N1226, N830);
xor XOR2 (N1245, N1243, N451);
buf BUF1 (N1246, N1234);
nor NOR4 (N1247, N1245, N1052, N443, N925);
and AND4 (N1248, N1246, N310, N815, N590);
or OR4 (N1249, N1218, N717, N452, N530);
xor XOR2 (N1250, N1239, N364);
nand NAND3 (N1251, N1237, N63, N524);
buf BUF1 (N1252, N1249);
buf BUF1 (N1253, N1252);
nor NOR3 (N1254, N1240, N1190, N1015);
nor NOR3 (N1255, N1250, N723, N151);
buf BUF1 (N1256, N1244);
and AND3 (N1257, N1256, N794, N1061);
xor XOR2 (N1258, N1228, N626);
and AND4 (N1259, N1257, N23, N183, N479);
nor NOR4 (N1260, N1251, N891, N922, N557);
nand NAND2 (N1261, N1258, N1067);
buf BUF1 (N1262, N1260);
buf BUF1 (N1263, N1242);
xor XOR2 (N1264, N1262, N241);
and AND3 (N1265, N1253, N453, N1169);
and AND2 (N1266, N1261, N1051);
and AND3 (N1267, N1264, N279, N773);
xor XOR2 (N1268, N1266, N744);
nand NAND3 (N1269, N1248, N213, N1189);
and AND2 (N1270, N1269, N938);
buf BUF1 (N1271, N1236);
or OR2 (N1272, N1254, N902);
nor NOR4 (N1273, N1247, N1167, N1269, N137);
nand NAND3 (N1274, N1268, N1198, N593);
and AND4 (N1275, N1265, N1214, N465, N788);
and AND4 (N1276, N1255, N94, N27, N118);
xor XOR2 (N1277, N1267, N507);
xor XOR2 (N1278, N1273, N1023);
or OR4 (N1279, N1259, N597, N1092, N738);
nor NOR4 (N1280, N1274, N134, N341, N941);
nor NOR3 (N1281, N1276, N26, N713);
nor NOR2 (N1282, N1277, N1269);
xor XOR2 (N1283, N1281, N1138);
not NOT1 (N1284, N1271);
xor XOR2 (N1285, N1278, N937);
buf BUF1 (N1286, N1272);
xor XOR2 (N1287, N1284, N144);
buf BUF1 (N1288, N1286);
xor XOR2 (N1289, N1263, N683);
xor XOR2 (N1290, N1283, N788);
nor NOR3 (N1291, N1285, N1234, N182);
nor NOR3 (N1292, N1291, N166, N221);
not NOT1 (N1293, N1292);
buf BUF1 (N1294, N1293);
or OR3 (N1295, N1282, N517, N588);
nand NAND2 (N1296, N1275, N486);
xor XOR2 (N1297, N1295, N557);
not NOT1 (N1298, N1280);
or OR4 (N1299, N1288, N207, N1259, N389);
and AND3 (N1300, N1289, N338, N762);
or OR4 (N1301, N1298, N123, N1238, N93);
not NOT1 (N1302, N1294);
buf BUF1 (N1303, N1290);
buf BUF1 (N1304, N1301);
not NOT1 (N1305, N1279);
nand NAND4 (N1306, N1303, N889, N801, N1180);
xor XOR2 (N1307, N1287, N70);
nand NAND2 (N1308, N1305, N1293);
xor XOR2 (N1309, N1308, N288);
nand NAND2 (N1310, N1309, N139);
buf BUF1 (N1311, N1296);
xor XOR2 (N1312, N1311, N353);
or OR3 (N1313, N1302, N652, N487);
xor XOR2 (N1314, N1304, N934);
or OR4 (N1315, N1312, N395, N727, N942);
xor XOR2 (N1316, N1313, N1099);
and AND4 (N1317, N1314, N954, N742, N859);
xor XOR2 (N1318, N1299, N269);
xor XOR2 (N1319, N1310, N202);
not NOT1 (N1320, N1270);
and AND3 (N1321, N1317, N660, N885);
nor NOR4 (N1322, N1319, N219, N725, N805);
buf BUF1 (N1323, N1300);
and AND3 (N1324, N1306, N324, N601);
and AND3 (N1325, N1318, N769, N937);
nand NAND2 (N1326, N1322, N808);
nand NAND4 (N1327, N1316, N62, N353, N304);
buf BUF1 (N1328, N1327);
nand NAND4 (N1329, N1326, N599, N740, N179);
buf BUF1 (N1330, N1307);
and AND3 (N1331, N1321, N1020, N740);
or OR3 (N1332, N1320, N444, N935);
buf BUF1 (N1333, N1325);
or OR3 (N1334, N1328, N117, N685);
and AND3 (N1335, N1332, N365, N229);
or OR4 (N1336, N1333, N1208, N567, N723);
buf BUF1 (N1337, N1323);
and AND2 (N1338, N1329, N1099);
or OR3 (N1339, N1324, N1304, N1224);
not NOT1 (N1340, N1315);
xor XOR2 (N1341, N1335, N651);
not NOT1 (N1342, N1340);
nor NOR2 (N1343, N1331, N866);
nor NOR3 (N1344, N1338, N1256, N1260);
not NOT1 (N1345, N1330);
or OR2 (N1346, N1334, N1127);
and AND2 (N1347, N1339, N584);
and AND2 (N1348, N1344, N667);
nand NAND4 (N1349, N1336, N728, N159, N1151);
or OR4 (N1350, N1348, N750, N156, N1169);
nand NAND2 (N1351, N1346, N890);
not NOT1 (N1352, N1345);
and AND3 (N1353, N1349, N621, N983);
or OR4 (N1354, N1352, N135, N299, N931);
nor NOR2 (N1355, N1342, N80);
nand NAND4 (N1356, N1337, N1167, N365, N191);
xor XOR2 (N1357, N1353, N517);
buf BUF1 (N1358, N1351);
or OR4 (N1359, N1341, N1049, N688, N579);
buf BUF1 (N1360, N1359);
and AND3 (N1361, N1354, N769, N654);
buf BUF1 (N1362, N1361);
xor XOR2 (N1363, N1357, N533);
buf BUF1 (N1364, N1360);
and AND3 (N1365, N1362, N1179, N431);
or OR4 (N1366, N1355, N215, N1074, N157);
or OR2 (N1367, N1297, N372);
not NOT1 (N1368, N1363);
xor XOR2 (N1369, N1365, N1266);
nand NAND4 (N1370, N1356, N494, N438, N513);
buf BUF1 (N1371, N1368);
nor NOR2 (N1372, N1366, N250);
or OR3 (N1373, N1372, N651, N120);
or OR2 (N1374, N1350, N96);
not NOT1 (N1375, N1367);
or OR2 (N1376, N1370, N912);
buf BUF1 (N1377, N1373);
buf BUF1 (N1378, N1347);
and AND2 (N1379, N1364, N46);
not NOT1 (N1380, N1377);
xor XOR2 (N1381, N1358, N971);
nand NAND3 (N1382, N1379, N652, N748);
nor NOR2 (N1383, N1380, N470);
nand NAND2 (N1384, N1382, N132);
xor XOR2 (N1385, N1383, N291);
nand NAND3 (N1386, N1369, N335, N186);
not NOT1 (N1387, N1374);
nor NOR2 (N1388, N1387, N140);
xor XOR2 (N1389, N1385, N502);
not NOT1 (N1390, N1384);
or OR3 (N1391, N1381, N956, N383);
and AND2 (N1392, N1390, N67);
nor NOR4 (N1393, N1371, N154, N282, N862);
and AND4 (N1394, N1391, N1207, N40, N1090);
not NOT1 (N1395, N1378);
or OR2 (N1396, N1343, N751);
xor XOR2 (N1397, N1394, N1360);
not NOT1 (N1398, N1397);
not NOT1 (N1399, N1396);
and AND4 (N1400, N1393, N278, N601, N1212);
nand NAND4 (N1401, N1388, N927, N469, N913);
and AND2 (N1402, N1400, N1391);
xor XOR2 (N1403, N1375, N983);
and AND2 (N1404, N1403, N335);
nand NAND3 (N1405, N1399, N961, N798);
xor XOR2 (N1406, N1398, N943);
nand NAND3 (N1407, N1389, N942, N320);
xor XOR2 (N1408, N1401, N455);
or OR4 (N1409, N1402, N242, N1237, N767);
nor NOR4 (N1410, N1405, N665, N636, N512);
xor XOR2 (N1411, N1392, N1081);
buf BUF1 (N1412, N1404);
xor XOR2 (N1413, N1412, N236);
not NOT1 (N1414, N1411);
xor XOR2 (N1415, N1409, N388);
or OR4 (N1416, N1410, N687, N1109, N551);
buf BUF1 (N1417, N1408);
not NOT1 (N1418, N1417);
nand NAND4 (N1419, N1414, N419, N1166, N1101);
nor NOR4 (N1420, N1407, N1025, N1097, N503);
and AND4 (N1421, N1419, N1327, N632, N538);
or OR4 (N1422, N1416, N676, N1381, N1395);
nand NAND4 (N1423, N349, N736, N892, N895);
buf BUF1 (N1424, N1406);
and AND2 (N1425, N1422, N1416);
buf BUF1 (N1426, N1386);
buf BUF1 (N1427, N1420);
and AND2 (N1428, N1415, N1427);
nand NAND2 (N1429, N948, N58);
or OR2 (N1430, N1418, N586);
and AND3 (N1431, N1428, N351, N5);
nand NAND4 (N1432, N1430, N503, N535, N580);
not NOT1 (N1433, N1424);
or OR3 (N1434, N1421, N786, N263);
and AND4 (N1435, N1423, N726, N798, N645);
and AND2 (N1436, N1426, N1363);
nand NAND4 (N1437, N1413, N211, N142, N926);
buf BUF1 (N1438, N1425);
and AND4 (N1439, N1437, N519, N247, N393);
nor NOR4 (N1440, N1431, N820, N372, N527);
or OR2 (N1441, N1432, N149);
and AND3 (N1442, N1438, N724, N72);
and AND3 (N1443, N1436, N313, N1030);
or OR2 (N1444, N1442, N983);
nand NAND3 (N1445, N1376, N1035, N1202);
xor XOR2 (N1446, N1429, N1373);
nor NOR3 (N1447, N1434, N989, N938);
buf BUF1 (N1448, N1443);
buf BUF1 (N1449, N1445);
xor XOR2 (N1450, N1448, N528);
buf BUF1 (N1451, N1435);
and AND3 (N1452, N1450, N1199, N683);
xor XOR2 (N1453, N1441, N439);
and AND2 (N1454, N1447, N694);
or OR3 (N1455, N1433, N1312, N1059);
nand NAND2 (N1456, N1454, N1350);
nand NAND2 (N1457, N1446, N726);
xor XOR2 (N1458, N1449, N1203);
not NOT1 (N1459, N1452);
buf BUF1 (N1460, N1459);
nor NOR4 (N1461, N1453, N1323, N1109, N679);
buf BUF1 (N1462, N1458);
buf BUF1 (N1463, N1460);
nand NAND2 (N1464, N1457, N506);
and AND3 (N1465, N1461, N100, N1414);
nand NAND3 (N1466, N1444, N1223, N235);
nor NOR2 (N1467, N1455, N990);
nor NOR3 (N1468, N1465, N434, N724);
xor XOR2 (N1469, N1456, N1414);
or OR3 (N1470, N1464, N1352, N101);
xor XOR2 (N1471, N1466, N788);
buf BUF1 (N1472, N1471);
nand NAND4 (N1473, N1469, N680, N1022, N1414);
nand NAND2 (N1474, N1463, N537);
xor XOR2 (N1475, N1474, N622);
buf BUF1 (N1476, N1473);
or OR3 (N1477, N1468, N174, N107);
or OR4 (N1478, N1451, N970, N521, N377);
nor NOR4 (N1479, N1477, N612, N1164, N1003);
or OR3 (N1480, N1476, N421, N594);
and AND3 (N1481, N1479, N969, N746);
nand NAND4 (N1482, N1470, N707, N599, N823);
or OR4 (N1483, N1482, N938, N297, N147);
not NOT1 (N1484, N1480);
and AND4 (N1485, N1462, N199, N228, N452);
nor NOR4 (N1486, N1467, N1375, N1427, N201);
nand NAND3 (N1487, N1484, N49, N876);
xor XOR2 (N1488, N1486, N420);
nor NOR2 (N1489, N1439, N965);
nand NAND2 (N1490, N1475, N821);
buf BUF1 (N1491, N1490);
and AND2 (N1492, N1485, N676);
buf BUF1 (N1493, N1440);
nand NAND3 (N1494, N1492, N429, N436);
or OR4 (N1495, N1493, N142, N1192, N1275);
xor XOR2 (N1496, N1487, N799);
not NOT1 (N1497, N1494);
or OR2 (N1498, N1488, N35);
and AND3 (N1499, N1483, N1238, N894);
nor NOR3 (N1500, N1481, N842, N1074);
buf BUF1 (N1501, N1499);
xor XOR2 (N1502, N1491, N1243);
buf BUF1 (N1503, N1472);
xor XOR2 (N1504, N1500, N86);
nor NOR4 (N1505, N1495, N1484, N1492, N920);
or OR3 (N1506, N1478, N878, N937);
nand NAND4 (N1507, N1503, N513, N745, N987);
nor NOR3 (N1508, N1505, N1166, N283);
not NOT1 (N1509, N1504);
nor NOR2 (N1510, N1508, N371);
xor XOR2 (N1511, N1496, N354);
nand NAND3 (N1512, N1511, N1483, N833);
or OR3 (N1513, N1512, N1093, N1369);
buf BUF1 (N1514, N1497);
buf BUF1 (N1515, N1498);
buf BUF1 (N1516, N1489);
not NOT1 (N1517, N1506);
buf BUF1 (N1518, N1502);
buf BUF1 (N1519, N1510);
not NOT1 (N1520, N1518);
nand NAND4 (N1521, N1501, N1122, N1437, N139);
xor XOR2 (N1522, N1513, N891);
not NOT1 (N1523, N1519);
xor XOR2 (N1524, N1520, N1166);
nor NOR3 (N1525, N1521, N66, N1185);
and AND4 (N1526, N1517, N317, N84, N46);
or OR2 (N1527, N1522, N1166);
xor XOR2 (N1528, N1516, N412);
and AND3 (N1529, N1528, N657, N381);
nor NOR3 (N1530, N1526, N440, N1331);
nand NAND4 (N1531, N1527, N312, N851, N178);
not NOT1 (N1532, N1530);
buf BUF1 (N1533, N1509);
and AND4 (N1534, N1525, N1460, N1102, N1191);
nor NOR3 (N1535, N1523, N1525, N736);
nor NOR3 (N1536, N1507, N265, N172);
not NOT1 (N1537, N1514);
and AND2 (N1538, N1529, N399);
nor NOR2 (N1539, N1534, N279);
or OR2 (N1540, N1537, N853);
nand NAND4 (N1541, N1538, N13, N1366, N434);
nor NOR4 (N1542, N1515, N1256, N1192, N1142);
nor NOR3 (N1543, N1536, N730, N656);
nand NAND3 (N1544, N1531, N1335, N815);
not NOT1 (N1545, N1543);
nor NOR2 (N1546, N1532, N34);
nand NAND3 (N1547, N1542, N262, N716);
nor NOR2 (N1548, N1547, N169);
not NOT1 (N1549, N1548);
xor XOR2 (N1550, N1544, N212);
nand NAND3 (N1551, N1541, N373, N1437);
xor XOR2 (N1552, N1545, N1075);
xor XOR2 (N1553, N1539, N1110);
nand NAND4 (N1554, N1533, N50, N359, N9);
not NOT1 (N1555, N1546);
xor XOR2 (N1556, N1553, N306);
not NOT1 (N1557, N1554);
buf BUF1 (N1558, N1524);
xor XOR2 (N1559, N1557, N451);
xor XOR2 (N1560, N1552, N1421);
or OR4 (N1561, N1556, N595, N572, N1096);
buf BUF1 (N1562, N1540);
and AND4 (N1563, N1559, N1003, N363, N101);
xor XOR2 (N1564, N1555, N553);
xor XOR2 (N1565, N1562, N696);
buf BUF1 (N1566, N1551);
nor NOR4 (N1567, N1560, N894, N1220, N1353);
not NOT1 (N1568, N1535);
and AND4 (N1569, N1550, N1098, N892, N1381);
buf BUF1 (N1570, N1567);
and AND3 (N1571, N1568, N648, N331);
nand NAND2 (N1572, N1558, N1492);
nand NAND4 (N1573, N1564, N532, N8, N1469);
buf BUF1 (N1574, N1549);
nor NOR3 (N1575, N1574, N694, N283);
nor NOR2 (N1576, N1570, N509);
nor NOR3 (N1577, N1571, N1463, N648);
nand NAND3 (N1578, N1576, N571, N218);
and AND3 (N1579, N1569, N397, N214);
and AND3 (N1580, N1561, N900, N689);
nand NAND2 (N1581, N1572, N1347);
nand NAND3 (N1582, N1577, N162, N1194);
buf BUF1 (N1583, N1578);
nor NOR3 (N1584, N1580, N399, N1564);
nand NAND3 (N1585, N1575, N803, N469);
or OR4 (N1586, N1583, N1311, N1385, N230);
or OR4 (N1587, N1563, N1301, N1178, N1339);
not NOT1 (N1588, N1573);
or OR3 (N1589, N1566, N58, N795);
and AND2 (N1590, N1589, N648);
and AND4 (N1591, N1585, N1077, N1571, N609);
not NOT1 (N1592, N1579);
xor XOR2 (N1593, N1588, N1289);
and AND2 (N1594, N1593, N1107);
nand NAND4 (N1595, N1581, N118, N548, N1377);
and AND3 (N1596, N1565, N1504, N413);
nor NOR2 (N1597, N1591, N486);
nand NAND4 (N1598, N1587, N1485, N356, N18);
nor NOR2 (N1599, N1586, N1593);
and AND3 (N1600, N1582, N742, N801);
nor NOR4 (N1601, N1598, N217, N1274, N156);
xor XOR2 (N1602, N1596, N1427);
xor XOR2 (N1603, N1590, N606);
buf BUF1 (N1604, N1601);
or OR4 (N1605, N1604, N400, N1078, N538);
xor XOR2 (N1606, N1592, N294);
xor XOR2 (N1607, N1600, N1078);
xor XOR2 (N1608, N1597, N637);
buf BUF1 (N1609, N1599);
buf BUF1 (N1610, N1608);
not NOT1 (N1611, N1606);
nand NAND3 (N1612, N1584, N158, N1345);
and AND3 (N1613, N1602, N806, N1474);
buf BUF1 (N1614, N1607);
buf BUF1 (N1615, N1613);
nand NAND3 (N1616, N1611, N1078, N1324);
buf BUF1 (N1617, N1595);
xor XOR2 (N1618, N1609, N1452);
and AND4 (N1619, N1612, N424, N1214, N1412);
nand NAND2 (N1620, N1617, N295);
and AND2 (N1621, N1620, N311);
not NOT1 (N1622, N1614);
and AND3 (N1623, N1610, N1439, N1361);
nand NAND4 (N1624, N1605, N1249, N1203, N361);
nand NAND2 (N1625, N1623, N393);
nor NOR3 (N1626, N1625, N1467, N1412);
not NOT1 (N1627, N1622);
not NOT1 (N1628, N1594);
and AND4 (N1629, N1618, N1388, N1604, N235);
nor NOR3 (N1630, N1627, N759, N233);
or OR4 (N1631, N1626, N682, N578, N1252);
not NOT1 (N1632, N1630);
xor XOR2 (N1633, N1619, N503);
or OR2 (N1634, N1633, N570);
and AND3 (N1635, N1629, N443, N135);
buf BUF1 (N1636, N1632);
nor NOR4 (N1637, N1624, N1393, N932, N773);
not NOT1 (N1638, N1631);
buf BUF1 (N1639, N1635);
and AND2 (N1640, N1616, N1180);
and AND2 (N1641, N1637, N1282);
not NOT1 (N1642, N1621);
not NOT1 (N1643, N1634);
not NOT1 (N1644, N1628);
buf BUF1 (N1645, N1636);
nor NOR3 (N1646, N1603, N576, N283);
xor XOR2 (N1647, N1642, N1152);
nor NOR3 (N1648, N1615, N1583, N188);
and AND2 (N1649, N1639, N602);
xor XOR2 (N1650, N1648, N1472);
and AND2 (N1651, N1649, N895);
nor NOR2 (N1652, N1644, N621);
not NOT1 (N1653, N1652);
nor NOR4 (N1654, N1645, N858, N1624, N337);
xor XOR2 (N1655, N1651, N419);
and AND4 (N1656, N1646, N1624, N1461, N269);
nand NAND3 (N1657, N1655, N847, N431);
or OR4 (N1658, N1656, N772, N948, N679);
not NOT1 (N1659, N1658);
nand NAND3 (N1660, N1654, N994, N1143);
or OR4 (N1661, N1640, N511, N793, N190);
nor NOR4 (N1662, N1660, N1387, N1461, N536);
and AND2 (N1663, N1641, N413);
or OR3 (N1664, N1643, N1309, N1083);
buf BUF1 (N1665, N1657);
nand NAND2 (N1666, N1650, N1535);
buf BUF1 (N1667, N1663);
and AND2 (N1668, N1666, N1087);
xor XOR2 (N1669, N1661, N1409);
nor NOR3 (N1670, N1659, N1440, N380);
not NOT1 (N1671, N1667);
xor XOR2 (N1672, N1669, N430);
nor NOR3 (N1673, N1672, N688, N544);
not NOT1 (N1674, N1671);
nand NAND3 (N1675, N1653, N714, N1239);
and AND2 (N1676, N1638, N1338);
nor NOR4 (N1677, N1662, N1467, N501, N1047);
xor XOR2 (N1678, N1676, N1671);
xor XOR2 (N1679, N1677, N418);
xor XOR2 (N1680, N1647, N1182);
not NOT1 (N1681, N1680);
not NOT1 (N1682, N1673);
and AND4 (N1683, N1670, N1377, N1633, N1620);
not NOT1 (N1684, N1679);
and AND3 (N1685, N1682, N1169, N224);
or OR2 (N1686, N1675, N1209);
or OR2 (N1687, N1674, N728);
or OR2 (N1688, N1668, N1491);
not NOT1 (N1689, N1684);
or OR4 (N1690, N1685, N596, N411, N339);
not NOT1 (N1691, N1681);
and AND3 (N1692, N1689, N1140, N395);
or OR2 (N1693, N1686, N671);
nor NOR4 (N1694, N1678, N177, N291, N889);
xor XOR2 (N1695, N1692, N276);
nor NOR2 (N1696, N1693, N1329);
nand NAND4 (N1697, N1687, N733, N582, N1175);
not NOT1 (N1698, N1688);
not NOT1 (N1699, N1665);
nor NOR4 (N1700, N1690, N416, N945, N210);
nand NAND4 (N1701, N1664, N108, N101, N758);
nor NOR4 (N1702, N1691, N645, N1413, N1183);
or OR3 (N1703, N1698, N804, N222);
buf BUF1 (N1704, N1699);
xor XOR2 (N1705, N1697, N545);
and AND4 (N1706, N1701, N1177, N306, N760);
buf BUF1 (N1707, N1705);
xor XOR2 (N1708, N1696, N1479);
nand NAND3 (N1709, N1683, N286, N199);
nor NOR2 (N1710, N1707, N725);
nor NOR2 (N1711, N1702, N874);
buf BUF1 (N1712, N1704);
buf BUF1 (N1713, N1709);
buf BUF1 (N1714, N1711);
nand NAND2 (N1715, N1712, N255);
xor XOR2 (N1716, N1700, N533);
buf BUF1 (N1717, N1713);
nor NOR4 (N1718, N1695, N868, N1262, N648);
buf BUF1 (N1719, N1710);
nand NAND3 (N1720, N1715, N58, N809);
buf BUF1 (N1721, N1708);
not NOT1 (N1722, N1719);
not NOT1 (N1723, N1714);
or OR4 (N1724, N1722, N508, N1544, N205);
buf BUF1 (N1725, N1718);
nor NOR2 (N1726, N1703, N530);
xor XOR2 (N1727, N1725, N841);
nor NOR3 (N1728, N1720, N262, N1147);
nor NOR2 (N1729, N1723, N961);
not NOT1 (N1730, N1721);
and AND3 (N1731, N1728, N353, N51);
and AND2 (N1732, N1729, N1520);
or OR4 (N1733, N1716, N1483, N429, N1014);
and AND3 (N1734, N1717, N1158, N1447);
xor XOR2 (N1735, N1706, N915);
xor XOR2 (N1736, N1726, N1121);
not NOT1 (N1737, N1731);
xor XOR2 (N1738, N1733, N1252);
and AND4 (N1739, N1727, N641, N1325, N379);
buf BUF1 (N1740, N1735);
xor XOR2 (N1741, N1694, N395);
not NOT1 (N1742, N1730);
buf BUF1 (N1743, N1739);
buf BUF1 (N1744, N1741);
nand NAND2 (N1745, N1734, N275);
buf BUF1 (N1746, N1737);
nor NOR2 (N1747, N1738, N31);
nand NAND2 (N1748, N1747, N824);
nand NAND3 (N1749, N1748, N1623, N921);
nand NAND4 (N1750, N1732, N1139, N264, N995);
nor NOR4 (N1751, N1742, N118, N703, N718);
xor XOR2 (N1752, N1744, N783);
and AND3 (N1753, N1724, N377, N631);
and AND2 (N1754, N1752, N921);
or OR2 (N1755, N1753, N1574);
or OR3 (N1756, N1751, N1493, N1743);
nor NOR2 (N1757, N1315, N1382);
xor XOR2 (N1758, N1749, N47);
nand NAND2 (N1759, N1745, N702);
buf BUF1 (N1760, N1754);
buf BUF1 (N1761, N1758);
not NOT1 (N1762, N1746);
buf BUF1 (N1763, N1757);
or OR4 (N1764, N1760, N445, N1052, N1200);
nand NAND4 (N1765, N1750, N164, N864, N1408);
nand NAND3 (N1766, N1736, N1596, N1213);
or OR3 (N1767, N1740, N1418, N1765);
nor NOR2 (N1768, N1549, N353);
and AND4 (N1769, N1755, N409, N66, N15);
xor XOR2 (N1770, N1767, N1590);
not NOT1 (N1771, N1764);
xor XOR2 (N1772, N1761, N263);
xor XOR2 (N1773, N1769, N104);
xor XOR2 (N1774, N1770, N1545);
nand NAND3 (N1775, N1766, N1648, N746);
nor NOR3 (N1776, N1772, N1287, N1712);
not NOT1 (N1777, N1768);
xor XOR2 (N1778, N1774, N1725);
nand NAND2 (N1779, N1763, N1739);
nor NOR3 (N1780, N1776, N769, N1624);
nor NOR4 (N1781, N1773, N1746, N1455, N1536);
not NOT1 (N1782, N1775);
and AND2 (N1783, N1781, N984);
and AND3 (N1784, N1759, N463, N1056);
or OR2 (N1785, N1778, N712);
or OR3 (N1786, N1780, N596, N1263);
nand NAND2 (N1787, N1786, N192);
not NOT1 (N1788, N1762);
nand NAND2 (N1789, N1777, N1155);
nor NOR2 (N1790, N1779, N129);
and AND3 (N1791, N1771, N36, N182);
nor NOR3 (N1792, N1788, N1281, N960);
not NOT1 (N1793, N1792);
and AND2 (N1794, N1791, N36);
nor NOR4 (N1795, N1782, N5, N1468, N337);
xor XOR2 (N1796, N1756, N81);
not NOT1 (N1797, N1795);
nor NOR3 (N1798, N1785, N809, N994);
nor NOR2 (N1799, N1790, N1222);
buf BUF1 (N1800, N1784);
or OR2 (N1801, N1787, N705);
buf BUF1 (N1802, N1793);
buf BUF1 (N1803, N1798);
nor NOR3 (N1804, N1800, N1132, N637);
buf BUF1 (N1805, N1783);
or OR2 (N1806, N1789, N1001);
nor NOR2 (N1807, N1803, N997);
nor NOR3 (N1808, N1799, N1261, N1083);
buf BUF1 (N1809, N1807);
buf BUF1 (N1810, N1806);
and AND4 (N1811, N1805, N1707, N326, N805);
or OR4 (N1812, N1796, N358, N938, N888);
nor NOR2 (N1813, N1810, N147);
and AND3 (N1814, N1801, N908, N1540);
nor NOR3 (N1815, N1812, N724, N281);
nor NOR2 (N1816, N1802, N1491);
not NOT1 (N1817, N1811);
not NOT1 (N1818, N1815);
or OR4 (N1819, N1814, N570, N186, N64);
nor NOR2 (N1820, N1818, N1724);
nand NAND3 (N1821, N1817, N220, N124);
xor XOR2 (N1822, N1794, N1598);
nand NAND3 (N1823, N1819, N1443, N1661);
xor XOR2 (N1824, N1809, N542);
buf BUF1 (N1825, N1808);
nand NAND4 (N1826, N1797, N74, N1425, N1323);
nand NAND4 (N1827, N1826, N1442, N1111, N850);
and AND4 (N1828, N1824, N1380, N1411, N731);
nor NOR3 (N1829, N1813, N1146, N1272);
or OR3 (N1830, N1816, N1252, N1113);
or OR4 (N1831, N1825, N950, N1322, N223);
and AND4 (N1832, N1804, N1613, N1302, N194);
buf BUF1 (N1833, N1830);
nand NAND4 (N1834, N1822, N1127, N1123, N206);
not NOT1 (N1835, N1829);
nor NOR4 (N1836, N1827, N931, N1832, N166);
and AND3 (N1837, N1803, N1799, N1086);
and AND3 (N1838, N1823, N1484, N365);
not NOT1 (N1839, N1837);
nor NOR3 (N1840, N1833, N1131, N1047);
xor XOR2 (N1841, N1839, N1448);
xor XOR2 (N1842, N1834, N990);
not NOT1 (N1843, N1838);
buf BUF1 (N1844, N1821);
or OR4 (N1845, N1843, N223, N952, N1680);
and AND4 (N1846, N1828, N1692, N1428, N665);
and AND4 (N1847, N1840, N257, N201, N617);
and AND3 (N1848, N1845, N1714, N686);
not NOT1 (N1849, N1820);
nor NOR4 (N1850, N1835, N1291, N512, N520);
nand NAND4 (N1851, N1846, N88, N701, N905);
buf BUF1 (N1852, N1844);
xor XOR2 (N1853, N1848, N1602);
nand NAND4 (N1854, N1847, N1694, N1574, N384);
nor NOR2 (N1855, N1854, N87);
or OR2 (N1856, N1855, N443);
xor XOR2 (N1857, N1831, N1117);
not NOT1 (N1858, N1851);
buf BUF1 (N1859, N1858);
not NOT1 (N1860, N1856);
not NOT1 (N1861, N1842);
nand NAND4 (N1862, N1836, N942, N173, N322);
xor XOR2 (N1863, N1849, N399);
nand NAND3 (N1864, N1862, N197, N96);
nor NOR2 (N1865, N1860, N1317);
and AND2 (N1866, N1864, N108);
xor XOR2 (N1867, N1865, N848);
nor NOR3 (N1868, N1853, N520, N962);
xor XOR2 (N1869, N1863, N1026);
not NOT1 (N1870, N1868);
or OR2 (N1871, N1869, N1304);
buf BUF1 (N1872, N1861);
nor NOR3 (N1873, N1857, N867, N835);
nor NOR4 (N1874, N1852, N74, N351, N303);
nand NAND3 (N1875, N1850, N910, N1470);
buf BUF1 (N1876, N1870);
buf BUF1 (N1877, N1874);
nand NAND4 (N1878, N1872, N1076, N1472, N1091);
or OR2 (N1879, N1871, N1534);
nand NAND3 (N1880, N1873, N1518, N943);
nor NOR3 (N1881, N1878, N713, N212);
nor NOR3 (N1882, N1866, N1265, N275);
nor NOR2 (N1883, N1859, N347);
and AND2 (N1884, N1877, N114);
xor XOR2 (N1885, N1841, N906);
nor NOR3 (N1886, N1879, N922, N25);
buf BUF1 (N1887, N1876);
nand NAND3 (N1888, N1867, N775, N1602);
and AND2 (N1889, N1886, N1258);
nand NAND3 (N1890, N1887, N1585, N939);
nand NAND4 (N1891, N1888, N1451, N156, N83);
and AND4 (N1892, N1891, N1652, N590, N351);
or OR3 (N1893, N1889, N362, N996);
nand NAND3 (N1894, N1880, N1497, N1595);
not NOT1 (N1895, N1893);
nor NOR2 (N1896, N1884, N1771);
xor XOR2 (N1897, N1881, N1729);
nor NOR4 (N1898, N1885, N1349, N650, N511);
buf BUF1 (N1899, N1892);
not NOT1 (N1900, N1896);
or OR4 (N1901, N1890, N255, N1276, N1716);
nand NAND4 (N1902, N1882, N418, N1450, N1050);
xor XOR2 (N1903, N1900, N1230);
buf BUF1 (N1904, N1903);
and AND3 (N1905, N1902, N989, N1836);
or OR2 (N1906, N1875, N490);
not NOT1 (N1907, N1906);
nor NOR4 (N1908, N1899, N966, N186, N1308);
buf BUF1 (N1909, N1894);
nand NAND2 (N1910, N1883, N46);
and AND2 (N1911, N1909, N1071);
nand NAND4 (N1912, N1910, N654, N735, N1033);
nand NAND4 (N1913, N1912, N1077, N856, N1621);
not NOT1 (N1914, N1907);
nor NOR4 (N1915, N1911, N83, N455, N1562);
nor NOR3 (N1916, N1898, N1813, N1119);
xor XOR2 (N1917, N1915, N1512);
nand NAND3 (N1918, N1904, N1889, N1034);
nand NAND3 (N1919, N1914, N242, N1849);
not NOT1 (N1920, N1918);
xor XOR2 (N1921, N1897, N1017);
nand NAND3 (N1922, N1908, N1406, N777);
nor NOR4 (N1923, N1917, N1800, N1603, N248);
not NOT1 (N1924, N1923);
nand NAND2 (N1925, N1919, N1434);
nand NAND3 (N1926, N1921, N761, N1739);
and AND2 (N1927, N1901, N1663);
buf BUF1 (N1928, N1913);
and AND2 (N1929, N1905, N1395);
nor NOR3 (N1930, N1928, N540, N1162);
nor NOR3 (N1931, N1916, N1199, N49);
nand NAND2 (N1932, N1922, N1898);
not NOT1 (N1933, N1920);
not NOT1 (N1934, N1932);
nor NOR2 (N1935, N1933, N985);
not NOT1 (N1936, N1935);
nand NAND3 (N1937, N1936, N1705, N190);
nand NAND2 (N1938, N1930, N1087);
not NOT1 (N1939, N1929);
and AND4 (N1940, N1925, N1936, N1578, N966);
not NOT1 (N1941, N1938);
xor XOR2 (N1942, N1927, N883);
not NOT1 (N1943, N1895);
xor XOR2 (N1944, N1940, N91);
and AND3 (N1945, N1941, N1618, N1138);
xor XOR2 (N1946, N1942, N85);
nand NAND4 (N1947, N1924, N85, N610, N885);
nor NOR2 (N1948, N1943, N727);
and AND4 (N1949, N1931, N1619, N805, N1488);
and AND2 (N1950, N1949, N538);
or OR4 (N1951, N1946, N1624, N1152, N1590);
buf BUF1 (N1952, N1939);
and AND4 (N1953, N1947, N764, N585, N1065);
or OR4 (N1954, N1944, N1409, N166, N687);
and AND4 (N1955, N1945, N158, N1800, N1859);
buf BUF1 (N1956, N1948);
nor NOR4 (N1957, N1956, N1027, N364, N1527);
or OR4 (N1958, N1957, N1266, N1573, N492);
xor XOR2 (N1959, N1958, N213);
nand NAND3 (N1960, N1950, N927, N817);
nor NOR4 (N1961, N1951, N664, N871, N1650);
buf BUF1 (N1962, N1953);
buf BUF1 (N1963, N1961);
nor NOR4 (N1964, N1963, N659, N830, N514);
nand NAND3 (N1965, N1952, N1607, N1517);
xor XOR2 (N1966, N1962, N1852);
and AND4 (N1967, N1959, N910, N1553, N124);
xor XOR2 (N1968, N1937, N1004);
or OR4 (N1969, N1964, N833, N495, N551);
buf BUF1 (N1970, N1960);
or OR4 (N1971, N1968, N1598, N436, N1806);
or OR3 (N1972, N1970, N874, N1205);
or OR4 (N1973, N1972, N1809, N320, N1112);
buf BUF1 (N1974, N1971);
xor XOR2 (N1975, N1955, N272);
xor XOR2 (N1976, N1969, N1105);
or OR2 (N1977, N1926, N453);
and AND3 (N1978, N1934, N1790, N220);
or OR4 (N1979, N1978, N1028, N557, N503);
nor NOR4 (N1980, N1966, N860, N1540, N1329);
buf BUF1 (N1981, N1967);
not NOT1 (N1982, N1981);
nor NOR2 (N1983, N1979, N1369);
nand NAND2 (N1984, N1980, N813);
and AND4 (N1985, N1954, N219, N1872, N1743);
not NOT1 (N1986, N1975);
not NOT1 (N1987, N1977);
nor NOR3 (N1988, N1976, N234, N698);
xor XOR2 (N1989, N1985, N1927);
buf BUF1 (N1990, N1983);
or OR2 (N1991, N1989, N20);
xor XOR2 (N1992, N1982, N869);
not NOT1 (N1993, N1984);
nor NOR3 (N1994, N1974, N7, N205);
or OR2 (N1995, N1988, N780);
nand NAND4 (N1996, N1990, N1039, N1166, N1325);
nor NOR4 (N1997, N1995, N46, N127, N549);
and AND3 (N1998, N1987, N419, N1910);
nand NAND2 (N1999, N1993, N326);
and AND2 (N2000, N1973, N353);
buf BUF1 (N2001, N1986);
or OR4 (N2002, N1992, N1383, N1757, N1868);
buf BUF1 (N2003, N1997);
buf BUF1 (N2004, N1991);
nand NAND2 (N2005, N2003, N144);
buf BUF1 (N2006, N2001);
xor XOR2 (N2007, N1994, N1184);
xor XOR2 (N2008, N1996, N284);
nor NOR4 (N2009, N1965, N1694, N672, N777);
buf BUF1 (N2010, N1998);
and AND4 (N2011, N2002, N151, N198, N1694);
nor NOR2 (N2012, N2010, N971);
or OR4 (N2013, N2004, N243, N1300, N1440);
not NOT1 (N2014, N2008);
buf BUF1 (N2015, N2013);
or OR2 (N2016, N2006, N211);
nand NAND2 (N2017, N2009, N1696);
or OR3 (N2018, N1999, N539, N1330);
xor XOR2 (N2019, N2011, N1473);
buf BUF1 (N2020, N2017);
or OR4 (N2021, N2012, N1895, N751, N1567);
xor XOR2 (N2022, N2015, N1962);
and AND3 (N2023, N2019, N920, N1156);
and AND2 (N2024, N2016, N1485);
xor XOR2 (N2025, N2007, N997);
nand NAND3 (N2026, N2005, N1934, N1325);
not NOT1 (N2027, N2023);
and AND2 (N2028, N2000, N163);
xor XOR2 (N2029, N2024, N1789);
nor NOR2 (N2030, N2027, N325);
or OR2 (N2031, N2014, N458);
buf BUF1 (N2032, N2031);
not NOT1 (N2033, N2021);
xor XOR2 (N2034, N2025, N325);
nor NOR3 (N2035, N2018, N904, N686);
not NOT1 (N2036, N2026);
buf BUF1 (N2037, N2020);
buf BUF1 (N2038, N2034);
nor NOR3 (N2039, N2033, N1169, N936);
nand NAND2 (N2040, N2028, N1191);
xor XOR2 (N2041, N2029, N1648);
and AND3 (N2042, N2037, N2016, N443);
not NOT1 (N2043, N2040);
nor NOR2 (N2044, N2039, N1516);
and AND4 (N2045, N2032, N60, N732, N1075);
nand NAND2 (N2046, N2045, N1379);
or OR2 (N2047, N2038, N1798);
and AND3 (N2048, N2035, N1947, N1151);
and AND3 (N2049, N2044, N1834, N694);
nor NOR2 (N2050, N2041, N347);
not NOT1 (N2051, N2048);
and AND2 (N2052, N2030, N975);
nor NOR2 (N2053, N2043, N1385);
and AND4 (N2054, N2022, N1586, N1772, N608);
nand NAND2 (N2055, N2052, N220);
xor XOR2 (N2056, N2050, N717);
xor XOR2 (N2057, N2042, N265);
nor NOR4 (N2058, N2053, N1750, N1939, N1134);
or OR2 (N2059, N2054, N1688);
not NOT1 (N2060, N2058);
xor XOR2 (N2061, N2046, N500);
buf BUF1 (N2062, N2051);
not NOT1 (N2063, N2059);
nor NOR2 (N2064, N2060, N1223);
xor XOR2 (N2065, N2057, N1781);
nand NAND4 (N2066, N2061, N1179, N499, N914);
not NOT1 (N2067, N2036);
nor NOR3 (N2068, N2067, N628, N315);
xor XOR2 (N2069, N2055, N334);
or OR3 (N2070, N2062, N850, N697);
nor NOR3 (N2071, N2056, N1494, N1470);
nor NOR2 (N2072, N2063, N1260);
nand NAND4 (N2073, N2066, N1846, N155, N1692);
nor NOR3 (N2074, N2072, N1997, N527);
and AND2 (N2075, N2074, N1169);
buf BUF1 (N2076, N2049);
not NOT1 (N2077, N2073);
not NOT1 (N2078, N2075);
or OR3 (N2079, N2064, N147, N1119);
buf BUF1 (N2080, N2070);
nand NAND3 (N2081, N2077, N1722, N1940);
or OR3 (N2082, N2081, N836, N1251);
nand NAND3 (N2083, N2071, N780, N1130);
and AND3 (N2084, N2079, N144, N1820);
and AND4 (N2085, N2084, N316, N1774, N1388);
nand NAND2 (N2086, N2068, N373);
buf BUF1 (N2087, N2078);
xor XOR2 (N2088, N2080, N1157);
xor XOR2 (N2089, N2069, N819);
nand NAND2 (N2090, N2047, N2016);
not NOT1 (N2091, N2076);
or OR4 (N2092, N2088, N845, N390, N1426);
nand NAND2 (N2093, N2082, N356);
nor NOR4 (N2094, N2083, N860, N1623, N1049);
not NOT1 (N2095, N2065);
or OR4 (N2096, N2090, N1986, N50, N937);
nor NOR4 (N2097, N2091, N40, N654, N1775);
buf BUF1 (N2098, N2096);
or OR3 (N2099, N2097, N1293, N917);
nor NOR4 (N2100, N2089, N1507, N534, N736);
or OR2 (N2101, N2100, N1856);
buf BUF1 (N2102, N2094);
nor NOR2 (N2103, N2087, N2035);
not NOT1 (N2104, N2086);
nor NOR4 (N2105, N2104, N756, N1158, N643);
not NOT1 (N2106, N2085);
or OR4 (N2107, N2098, N257, N1858, N1152);
and AND3 (N2108, N2107, N1769, N150);
or OR4 (N2109, N2103, N320, N1799, N1490);
not NOT1 (N2110, N2106);
and AND2 (N2111, N2092, N547);
and AND2 (N2112, N2093, N694);
and AND4 (N2113, N2102, N1886, N413, N390);
xor XOR2 (N2114, N2095, N1322);
and AND2 (N2115, N2110, N1523);
nor NOR4 (N2116, N2113, N15, N1921, N1658);
and AND3 (N2117, N2111, N571, N543);
nand NAND2 (N2118, N2117, N836);
or OR4 (N2119, N2108, N151, N481, N500);
nand NAND2 (N2120, N2099, N871);
buf BUF1 (N2121, N2116);
or OR4 (N2122, N2101, N1268, N1961, N881);
nor NOR4 (N2123, N2121, N1374, N624, N85);
or OR4 (N2124, N2115, N576, N1351, N1343);
nand NAND3 (N2125, N2112, N2030, N68);
and AND4 (N2126, N2105, N1689, N1553, N1264);
not NOT1 (N2127, N2124);
nor NOR4 (N2128, N2127, N600, N255, N885);
nor NOR4 (N2129, N2122, N1355, N1331, N902);
and AND4 (N2130, N2109, N1966, N1577, N1457);
and AND2 (N2131, N2128, N1859);
not NOT1 (N2132, N2129);
or OR4 (N2133, N2126, N260, N2103, N669);
not NOT1 (N2134, N2119);
buf BUF1 (N2135, N2114);
nor NOR4 (N2136, N2133, N2069, N1769, N1065);
buf BUF1 (N2137, N2135);
nand NAND3 (N2138, N2137, N627, N1756);
not NOT1 (N2139, N2120);
not NOT1 (N2140, N2134);
not NOT1 (N2141, N2132);
xor XOR2 (N2142, N2131, N600);
nor NOR2 (N2143, N2136, N531);
xor XOR2 (N2144, N2142, N1016);
buf BUF1 (N2145, N2118);
or OR3 (N2146, N2130, N2095, N1451);
buf BUF1 (N2147, N2144);
buf BUF1 (N2148, N2145);
or OR2 (N2149, N2123, N284);
xor XOR2 (N2150, N2141, N736);
nor NOR3 (N2151, N2147, N685, N248);
xor XOR2 (N2152, N2151, N1368);
nor NOR4 (N2153, N2139, N212, N1661, N1789);
not NOT1 (N2154, N2138);
xor XOR2 (N2155, N2153, N705);
and AND2 (N2156, N2143, N1849);
xor XOR2 (N2157, N2146, N1734);
or OR2 (N2158, N2150, N667);
nor NOR3 (N2159, N2155, N1988, N2088);
xor XOR2 (N2160, N2125, N474);
buf BUF1 (N2161, N2159);
or OR4 (N2162, N2140, N1803, N2142, N436);
nand NAND2 (N2163, N2156, N797);
nor NOR3 (N2164, N2158, N243, N1417);
and AND3 (N2165, N2163, N829, N915);
not NOT1 (N2166, N2161);
nor NOR3 (N2167, N2152, N1833, N1054);
or OR3 (N2168, N2160, N353, N1347);
not NOT1 (N2169, N2148);
nor NOR2 (N2170, N2162, N1713);
not NOT1 (N2171, N2157);
nand NAND3 (N2172, N2168, N1323, N1255);
nor NOR2 (N2173, N2166, N1318);
nor NOR4 (N2174, N2171, N1265, N1970, N1262);
not NOT1 (N2175, N2172);
nand NAND3 (N2176, N2149, N972, N1949);
nor NOR2 (N2177, N2167, N737);
buf BUF1 (N2178, N2173);
buf BUF1 (N2179, N2169);
not NOT1 (N2180, N2176);
buf BUF1 (N2181, N2164);
and AND2 (N2182, N2181, N825);
xor XOR2 (N2183, N2177, N2060);
nand NAND3 (N2184, N2179, N761, N1711);
nor NOR3 (N2185, N2154, N334, N1176);
xor XOR2 (N2186, N2183, N1929);
buf BUF1 (N2187, N2184);
nand NAND2 (N2188, N2180, N644);
and AND2 (N2189, N2175, N651);
nand NAND3 (N2190, N2186, N1025, N157);
or OR2 (N2191, N2174, N985);
nand NAND2 (N2192, N2191, N862);
nand NAND3 (N2193, N2188, N1084, N376);
not NOT1 (N2194, N2193);
not NOT1 (N2195, N2189);
xor XOR2 (N2196, N2195, N1738);
xor XOR2 (N2197, N2190, N1243);
nand NAND2 (N2198, N2196, N37);
buf BUF1 (N2199, N2165);
nor NOR3 (N2200, N2197, N1505, N2050);
or OR3 (N2201, N2178, N1020, N1628);
or OR4 (N2202, N2198, N848, N1584, N554);
and AND3 (N2203, N2202, N2126, N1018);
or OR4 (N2204, N2170, N1547, N466, N1931);
or OR4 (N2205, N2204, N389, N683, N1316);
and AND4 (N2206, N2205, N829, N2184, N358);
not NOT1 (N2207, N2187);
and AND4 (N2208, N2200, N531, N1597, N625);
nor NOR4 (N2209, N2206, N1325, N1193, N1703);
and AND3 (N2210, N2199, N2143, N85);
nor NOR3 (N2211, N2207, N1095, N1470);
xor XOR2 (N2212, N2203, N817);
xor XOR2 (N2213, N2182, N1387);
buf BUF1 (N2214, N2213);
nor NOR4 (N2215, N2192, N1143, N1142, N1533);
buf BUF1 (N2216, N2194);
or OR2 (N2217, N2209, N429);
xor XOR2 (N2218, N2217, N768);
not NOT1 (N2219, N2215);
not NOT1 (N2220, N2212);
buf BUF1 (N2221, N2201);
xor XOR2 (N2222, N2211, N1190);
nand NAND3 (N2223, N2185, N2114, N706);
or OR2 (N2224, N2214, N1416);
and AND4 (N2225, N2216, N2124, N1195, N540);
buf BUF1 (N2226, N2223);
or OR3 (N2227, N2224, N1121, N231);
buf BUF1 (N2228, N2210);
buf BUF1 (N2229, N2219);
or OR2 (N2230, N2229, N826);
nand NAND2 (N2231, N2225, N1117);
and AND2 (N2232, N2226, N1123);
nor NOR4 (N2233, N2232, N823, N1606, N697);
xor XOR2 (N2234, N2228, N1164);
buf BUF1 (N2235, N2222);
buf BUF1 (N2236, N2230);
nand NAND3 (N2237, N2221, N1546, N1968);
and AND4 (N2238, N2233, N1718, N1290, N1196);
buf BUF1 (N2239, N2227);
nor NOR4 (N2240, N2218, N1370, N1121, N9);
buf BUF1 (N2241, N2238);
nand NAND2 (N2242, N2239, N1589);
and AND2 (N2243, N2236, N1953);
xor XOR2 (N2244, N2231, N2007);
xor XOR2 (N2245, N2237, N1461);
xor XOR2 (N2246, N2245, N1896);
xor XOR2 (N2247, N2220, N1612);
nand NAND3 (N2248, N2244, N608, N734);
and AND2 (N2249, N2234, N1274);
or OR4 (N2250, N2241, N324, N149, N279);
nand NAND4 (N2251, N2208, N1307, N582, N1038);
or OR4 (N2252, N2246, N386, N1155, N1485);
xor XOR2 (N2253, N2250, N821);
nand NAND4 (N2254, N2247, N1346, N325, N583);
buf BUF1 (N2255, N2253);
nor NOR2 (N2256, N2254, N1172);
nand NAND2 (N2257, N2242, N684);
not NOT1 (N2258, N2240);
or OR3 (N2259, N2235, N283, N1512);
nor NOR4 (N2260, N2257, N320, N1253, N607);
nand NAND3 (N2261, N2258, N750, N1269);
nor NOR4 (N2262, N2243, N1842, N1692, N669);
not NOT1 (N2263, N2252);
and AND4 (N2264, N2262, N472, N1911, N282);
nor NOR4 (N2265, N2249, N2181, N1693, N1660);
or OR2 (N2266, N2251, N1578);
nand NAND3 (N2267, N2259, N2019, N1676);
nand NAND3 (N2268, N2248, N2195, N1417);
xor XOR2 (N2269, N2255, N153);
nand NAND3 (N2270, N2265, N269, N1355);
xor XOR2 (N2271, N2268, N2032);
buf BUF1 (N2272, N2263);
buf BUF1 (N2273, N2267);
not NOT1 (N2274, N2261);
xor XOR2 (N2275, N2274, N2164);
and AND3 (N2276, N2269, N1468, N1459);
not NOT1 (N2277, N2276);
xor XOR2 (N2278, N2264, N312);
xor XOR2 (N2279, N2275, N1587);
not NOT1 (N2280, N2271);
buf BUF1 (N2281, N2256);
xor XOR2 (N2282, N2270, N957);
nor NOR2 (N2283, N2260, N1130);
buf BUF1 (N2284, N2280);
buf BUF1 (N2285, N2279);
and AND3 (N2286, N2272, N1667, N120);
nor NOR4 (N2287, N2285, N1132, N1135, N1645);
and AND4 (N2288, N2284, N521, N1980, N158);
not NOT1 (N2289, N2273);
buf BUF1 (N2290, N2286);
or OR4 (N2291, N2289, N526, N1111, N1229);
xor XOR2 (N2292, N2287, N827);
and AND2 (N2293, N2282, N2136);
or OR2 (N2294, N2290, N1088);
nor NOR4 (N2295, N2277, N1307, N1005, N907);
xor XOR2 (N2296, N2281, N666);
nor NOR4 (N2297, N2266, N767, N726, N2158);
nor NOR4 (N2298, N2296, N796, N1873, N368);
xor XOR2 (N2299, N2291, N964);
nor NOR2 (N2300, N2298, N1459);
nand NAND2 (N2301, N2278, N237);
and AND2 (N2302, N2288, N1682);
not NOT1 (N2303, N2295);
or OR4 (N2304, N2299, N942, N1456, N72);
and AND2 (N2305, N2303, N1588);
and AND2 (N2306, N2305, N1851);
xor XOR2 (N2307, N2283, N1413);
nor NOR4 (N2308, N2304, N1408, N1081, N1364);
xor XOR2 (N2309, N2306, N222);
xor XOR2 (N2310, N2300, N223);
nor NOR4 (N2311, N2302, N775, N1981, N2264);
and AND3 (N2312, N2301, N78, N2000);
buf BUF1 (N2313, N2297);
nor NOR4 (N2314, N2292, N2117, N6, N267);
and AND2 (N2315, N2307, N627);
nor NOR3 (N2316, N2293, N2117, N2234);
or OR4 (N2317, N2314, N2245, N1362, N114);
or OR3 (N2318, N2317, N2028, N527);
nand NAND4 (N2319, N2310, N316, N926, N575);
buf BUF1 (N2320, N2315);
or OR4 (N2321, N2319, N234, N429, N936);
nor NOR2 (N2322, N2316, N2041);
and AND4 (N2323, N2308, N481, N1648, N1553);
not NOT1 (N2324, N2320);
xor XOR2 (N2325, N2313, N238);
xor XOR2 (N2326, N2324, N598);
nand NAND3 (N2327, N2323, N856, N1081);
or OR3 (N2328, N2321, N945, N418);
nand NAND3 (N2329, N2325, N2070, N2141);
nor NOR4 (N2330, N2322, N510, N2110, N1472);
buf BUF1 (N2331, N2318);
not NOT1 (N2332, N2311);
or OR3 (N2333, N2327, N954, N2209);
and AND2 (N2334, N2332, N170);
buf BUF1 (N2335, N2309);
and AND2 (N2336, N2294, N1851);
not NOT1 (N2337, N2329);
nor NOR2 (N2338, N2335, N995);
or OR2 (N2339, N2334, N380);
not NOT1 (N2340, N2312);
buf BUF1 (N2341, N2333);
nor NOR3 (N2342, N2336, N290, N1133);
and AND2 (N2343, N2342, N183);
xor XOR2 (N2344, N2328, N1900);
nor NOR3 (N2345, N2343, N991, N1148);
and AND4 (N2346, N2326, N2132, N1686, N1278);
not NOT1 (N2347, N2346);
nor NOR4 (N2348, N2341, N707, N876, N2346);
and AND3 (N2349, N2331, N1782, N584);
nor NOR4 (N2350, N2347, N1164, N108, N1308);
nor NOR3 (N2351, N2350, N297, N1417);
or OR3 (N2352, N2330, N199, N1367);
buf BUF1 (N2353, N2351);
xor XOR2 (N2354, N2352, N537);
nor NOR4 (N2355, N2340, N241, N2109, N2097);
buf BUF1 (N2356, N2353);
xor XOR2 (N2357, N2339, N1808);
nand NAND4 (N2358, N2345, N2017, N862, N528);
xor XOR2 (N2359, N2358, N2267);
or OR2 (N2360, N2348, N1429);
nand NAND2 (N2361, N2357, N1344);
and AND2 (N2362, N2355, N2246);
buf BUF1 (N2363, N2359);
xor XOR2 (N2364, N2344, N170);
nand NAND4 (N2365, N2356, N1682, N2118, N1261);
nand NAND2 (N2366, N2361, N933);
not NOT1 (N2367, N2364);
or OR3 (N2368, N2363, N1695, N17);
or OR4 (N2369, N2362, N1755, N1451, N862);
nand NAND3 (N2370, N2368, N547, N1923);
not NOT1 (N2371, N2369);
and AND2 (N2372, N2338, N775);
and AND3 (N2373, N2360, N682, N538);
or OR3 (N2374, N2366, N1295, N341);
nand NAND4 (N2375, N2373, N1362, N1240, N1495);
buf BUF1 (N2376, N2372);
xor XOR2 (N2377, N2349, N400);
not NOT1 (N2378, N2367);
nand NAND2 (N2379, N2371, N166);
and AND2 (N2380, N2377, N62);
and AND3 (N2381, N2379, N1611, N1167);
buf BUF1 (N2382, N2375);
nand NAND2 (N2383, N2365, N1289);
not NOT1 (N2384, N2381);
not NOT1 (N2385, N2370);
buf BUF1 (N2386, N2376);
buf BUF1 (N2387, N2382);
xor XOR2 (N2388, N2385, N661);
buf BUF1 (N2389, N2378);
xor XOR2 (N2390, N2384, N2105);
nor NOR4 (N2391, N2390, N1778, N1335, N959);
not NOT1 (N2392, N2388);
buf BUF1 (N2393, N2337);
nand NAND4 (N2394, N2386, N227, N1854, N2380);
not NOT1 (N2395, N1962);
or OR2 (N2396, N2389, N727);
nand NAND3 (N2397, N2383, N1953, N2125);
nand NAND4 (N2398, N2397, N1997, N523, N1068);
nor NOR2 (N2399, N2392, N2266);
or OR2 (N2400, N2374, N846);
xor XOR2 (N2401, N2395, N450);
and AND4 (N2402, N2391, N131, N503, N1259);
nor NOR2 (N2403, N2398, N1347);
xor XOR2 (N2404, N2393, N1074);
buf BUF1 (N2405, N2394);
or OR4 (N2406, N2401, N1055, N271, N679);
xor XOR2 (N2407, N2399, N1953);
xor XOR2 (N2408, N2407, N73);
or OR3 (N2409, N2387, N1411, N1597);
nor NOR4 (N2410, N2354, N1446, N575, N2340);
and AND2 (N2411, N2396, N341);
or OR4 (N2412, N2402, N1289, N201, N464);
nor NOR3 (N2413, N2406, N600, N823);
nand NAND2 (N2414, N2411, N1016);
nor NOR2 (N2415, N2414, N585);
and AND3 (N2416, N2405, N1697, N1403);
xor XOR2 (N2417, N2413, N81);
xor XOR2 (N2418, N2415, N653);
not NOT1 (N2419, N2409);
and AND3 (N2420, N2419, N1978, N1084);
nand NAND3 (N2421, N2418, N687, N765);
buf BUF1 (N2422, N2421);
nor NOR3 (N2423, N2412, N776, N1568);
or OR4 (N2424, N2423, N167, N977, N641);
xor XOR2 (N2425, N2400, N1292);
nor NOR4 (N2426, N2403, N174, N1094, N1395);
or OR2 (N2427, N2422, N1330);
or OR3 (N2428, N2408, N1036, N2198);
buf BUF1 (N2429, N2427);
nand NAND3 (N2430, N2426, N268, N1528);
not NOT1 (N2431, N2425);
xor XOR2 (N2432, N2431, N1530);
nand NAND4 (N2433, N2429, N1547, N686, N1219);
nand NAND2 (N2434, N2433, N1729);
xor XOR2 (N2435, N2410, N1190);
nor NOR4 (N2436, N2430, N11, N1033, N1672);
and AND2 (N2437, N2432, N772);
not NOT1 (N2438, N2437);
and AND2 (N2439, N2435, N1577);
buf BUF1 (N2440, N2404);
xor XOR2 (N2441, N2434, N1410);
and AND2 (N2442, N2424, N505);
or OR4 (N2443, N2439, N1614, N1395, N406);
nand NAND2 (N2444, N2428, N1323);
nor NOR3 (N2445, N2417, N2185, N1398);
nand NAND4 (N2446, N2443, N1726, N1205, N2336);
not NOT1 (N2447, N2444);
buf BUF1 (N2448, N2441);
not NOT1 (N2449, N2448);
nor NOR2 (N2450, N2436, N1973);
not NOT1 (N2451, N2450);
nor NOR3 (N2452, N2451, N246, N12);
not NOT1 (N2453, N2447);
not NOT1 (N2454, N2449);
buf BUF1 (N2455, N2445);
not NOT1 (N2456, N2438);
and AND4 (N2457, N2440, N1301, N757, N1333);
xor XOR2 (N2458, N2455, N685);
nand NAND3 (N2459, N2458, N2433, N580);
not NOT1 (N2460, N2456);
buf BUF1 (N2461, N2446);
or OR3 (N2462, N2460, N569, N288);
nand NAND3 (N2463, N2416, N432, N622);
nor NOR2 (N2464, N2463, N767);
and AND3 (N2465, N2457, N1669, N1270);
xor XOR2 (N2466, N2461, N961);
or OR4 (N2467, N2442, N1582, N177, N1492);
not NOT1 (N2468, N2462);
and AND2 (N2469, N2454, N446);
xor XOR2 (N2470, N2453, N1944);
and AND3 (N2471, N2467, N1755, N2129);
and AND3 (N2472, N2464, N774, N899);
or OR3 (N2473, N2465, N1860, N663);
nand NAND3 (N2474, N2466, N1248, N1781);
not NOT1 (N2475, N2452);
and AND3 (N2476, N2475, N2067, N1728);
xor XOR2 (N2477, N2469, N1709);
or OR3 (N2478, N2476, N29, N457);
buf BUF1 (N2479, N2468);
and AND3 (N2480, N2479, N5, N2320);
and AND2 (N2481, N2473, N1847);
nor NOR2 (N2482, N2471, N1450);
nand NAND4 (N2483, N2480, N1782, N476, N2321);
or OR2 (N2484, N2459, N1021);
xor XOR2 (N2485, N2472, N545);
buf BUF1 (N2486, N2485);
or OR2 (N2487, N2481, N1283);
and AND4 (N2488, N2487, N1266, N1686, N1013);
buf BUF1 (N2489, N2484);
not NOT1 (N2490, N2474);
buf BUF1 (N2491, N2477);
nor NOR2 (N2492, N2489, N999);
not NOT1 (N2493, N2420);
nand NAND4 (N2494, N2483, N826, N936, N788);
buf BUF1 (N2495, N2470);
nand NAND4 (N2496, N2494, N2381, N1577, N1958);
or OR4 (N2497, N2478, N837, N297, N919);
or OR2 (N2498, N2497, N275);
nor NOR2 (N2499, N2486, N1945);
not NOT1 (N2500, N2490);
nor NOR4 (N2501, N2495, N1409, N1465, N1034);
or OR4 (N2502, N2499, N727, N1834, N1823);
not NOT1 (N2503, N2501);
nand NAND4 (N2504, N2492, N1381, N1409, N1582);
and AND3 (N2505, N2491, N524, N1182);
xor XOR2 (N2506, N2482, N1981);
and AND2 (N2507, N2493, N1212);
buf BUF1 (N2508, N2504);
not NOT1 (N2509, N2488);
or OR4 (N2510, N2509, N812, N2113, N372);
xor XOR2 (N2511, N2510, N1181);
not NOT1 (N2512, N2508);
buf BUF1 (N2513, N2503);
nor NOR4 (N2514, N2513, N466, N2359, N1706);
nand NAND2 (N2515, N2511, N83);
nor NOR3 (N2516, N2500, N1718, N1521);
xor XOR2 (N2517, N2498, N194);
not NOT1 (N2518, N2517);
xor XOR2 (N2519, N2516, N1847);
or OR3 (N2520, N2505, N638, N560);
or OR2 (N2521, N2518, N2148);
nand NAND3 (N2522, N2502, N1208, N921);
nor NOR3 (N2523, N2496, N1169, N1916);
nand NAND2 (N2524, N2506, N243);
and AND2 (N2525, N2520, N2175);
buf BUF1 (N2526, N2523);
not NOT1 (N2527, N2524);
and AND2 (N2528, N2519, N232);
nor NOR4 (N2529, N2512, N1669, N95, N1747);
not NOT1 (N2530, N2525);
nor NOR4 (N2531, N2507, N1522, N1203, N998);
nand NAND2 (N2532, N2522, N515);
nor NOR3 (N2533, N2521, N965, N1085);
xor XOR2 (N2534, N2533, N1806);
and AND2 (N2535, N2529, N2077);
buf BUF1 (N2536, N2531);
and AND3 (N2537, N2528, N2408, N1676);
xor XOR2 (N2538, N2532, N1968);
and AND4 (N2539, N2527, N2165, N1335, N1776);
nand NAND3 (N2540, N2534, N547, N374);
not NOT1 (N2541, N2514);
not NOT1 (N2542, N2537);
nor NOR4 (N2543, N2542, N1313, N2224, N963);
xor XOR2 (N2544, N2539, N2186);
not NOT1 (N2545, N2536);
xor XOR2 (N2546, N2538, N1899);
nand NAND4 (N2547, N2515, N1964, N940, N1931);
or OR2 (N2548, N2530, N590);
nor NOR3 (N2549, N2526, N1626, N1365);
nand NAND2 (N2550, N2545, N720);
xor XOR2 (N2551, N2541, N1321);
not NOT1 (N2552, N2551);
not NOT1 (N2553, N2549);
nand NAND2 (N2554, N2544, N262);
and AND4 (N2555, N2554, N1288, N1557, N1585);
nor NOR4 (N2556, N2535, N1591, N970, N628);
not NOT1 (N2557, N2547);
nor NOR4 (N2558, N2553, N358, N1400, N519);
and AND4 (N2559, N2552, N1411, N957, N1086);
not NOT1 (N2560, N2540);
and AND3 (N2561, N2559, N1722, N215);
nand NAND3 (N2562, N2543, N2, N1554);
or OR4 (N2563, N2556, N2285, N2419, N260);
not NOT1 (N2564, N2562);
not NOT1 (N2565, N2546);
or OR2 (N2566, N2561, N1485);
and AND4 (N2567, N2548, N775, N2045, N2303);
buf BUF1 (N2568, N2563);
buf BUF1 (N2569, N2567);
xor XOR2 (N2570, N2564, N1896);
nor NOR3 (N2571, N2557, N1351, N260);
nor NOR4 (N2572, N2565, N568, N825, N237);
not NOT1 (N2573, N2568);
not NOT1 (N2574, N2569);
and AND3 (N2575, N2558, N2030, N2286);
and AND3 (N2576, N2555, N980, N401);
buf BUF1 (N2577, N2575);
nand NAND2 (N2578, N2550, N1524);
nor NOR2 (N2579, N2572, N2375);
and AND4 (N2580, N2570, N1029, N929, N2372);
xor XOR2 (N2581, N2578, N1746);
nor NOR3 (N2582, N2573, N2532, N1116);
or OR3 (N2583, N2577, N231, N1706);
or OR2 (N2584, N2560, N1628);
or OR4 (N2585, N2576, N290, N502, N994);
buf BUF1 (N2586, N2566);
nor NOR2 (N2587, N2579, N142);
nand NAND4 (N2588, N2574, N1343, N436, N587);
buf BUF1 (N2589, N2584);
xor XOR2 (N2590, N2571, N1419);
xor XOR2 (N2591, N2583, N974);
not NOT1 (N2592, N2581);
or OR4 (N2593, N2587, N2522, N1993, N1732);
buf BUF1 (N2594, N2592);
nand NAND2 (N2595, N2591, N1634);
buf BUF1 (N2596, N2585);
buf BUF1 (N2597, N2588);
nand NAND3 (N2598, N2593, N326, N1495);
nor NOR2 (N2599, N2597, N959);
xor XOR2 (N2600, N2595, N1200);
buf BUF1 (N2601, N2600);
and AND3 (N2602, N2601, N340, N2383);
buf BUF1 (N2603, N2594);
and AND3 (N2604, N2598, N192, N1372);
xor XOR2 (N2605, N2590, N1889);
and AND3 (N2606, N2589, N547, N1840);
nor NOR2 (N2607, N2604, N1243);
xor XOR2 (N2608, N2603, N1438);
and AND4 (N2609, N2586, N2433, N610, N619);
and AND3 (N2610, N2607, N2579, N985);
buf BUF1 (N2611, N2610);
buf BUF1 (N2612, N2602);
buf BUF1 (N2613, N2611);
buf BUF1 (N2614, N2606);
not NOT1 (N2615, N2609);
or OR4 (N2616, N2580, N1646, N1320, N2006);
nand NAND2 (N2617, N2613, N2046);
nand NAND3 (N2618, N2608, N2070, N1914);
nor NOR3 (N2619, N2614, N2586, N2552);
not NOT1 (N2620, N2582);
xor XOR2 (N2621, N2620, N1244);
xor XOR2 (N2622, N2617, N2509);
and AND4 (N2623, N2618, N1682, N1133, N1092);
or OR4 (N2624, N2605, N820, N1901, N373);
or OR4 (N2625, N2596, N2607, N218, N2410);
nand NAND2 (N2626, N2599, N1974);
nand NAND4 (N2627, N2624, N1160, N506, N75);
buf BUF1 (N2628, N2616);
and AND3 (N2629, N2626, N930, N2398);
nor NOR4 (N2630, N2622, N837, N2249, N283);
or OR2 (N2631, N2623, N1238);
xor XOR2 (N2632, N2612, N448);
nor NOR3 (N2633, N2632, N164, N2518);
nand NAND4 (N2634, N2615, N2400, N440, N69);
and AND4 (N2635, N2633, N2055, N1122, N1506);
nor NOR4 (N2636, N2621, N2108, N45, N260);
xor XOR2 (N2637, N2629, N1008);
nand NAND3 (N2638, N2631, N1711, N17);
xor XOR2 (N2639, N2636, N653);
or OR2 (N2640, N2635, N2600);
buf BUF1 (N2641, N2640);
xor XOR2 (N2642, N2619, N2155);
buf BUF1 (N2643, N2627);
nand NAND3 (N2644, N2639, N2581, N576);
buf BUF1 (N2645, N2643);
or OR2 (N2646, N2628, N1508);
or OR3 (N2647, N2642, N1122, N1109);
nor NOR3 (N2648, N2646, N599, N1245);
not NOT1 (N2649, N2630);
not NOT1 (N2650, N2647);
or OR4 (N2651, N2649, N197, N2309, N2630);
nand NAND3 (N2652, N2637, N130, N2606);
nand NAND3 (N2653, N2638, N1967, N1856);
nor NOR2 (N2654, N2645, N168);
buf BUF1 (N2655, N2644);
and AND2 (N2656, N2655, N2181);
nor NOR4 (N2657, N2650, N456, N2579, N1783);
nand NAND4 (N2658, N2653, N1523, N1431, N805);
nor NOR3 (N2659, N2641, N1052, N1771);
not NOT1 (N2660, N2651);
or OR3 (N2661, N2652, N1977, N47);
buf BUF1 (N2662, N2654);
or OR4 (N2663, N2634, N584, N334, N754);
xor XOR2 (N2664, N2657, N604);
and AND3 (N2665, N2648, N2100, N2310);
not NOT1 (N2666, N2659);
xor XOR2 (N2667, N2656, N1417);
not NOT1 (N2668, N2660);
not NOT1 (N2669, N2663);
or OR4 (N2670, N2661, N2191, N1241, N2430);
nand NAND2 (N2671, N2664, N160);
or OR4 (N2672, N2665, N2525, N1683, N2238);
nor NOR2 (N2673, N2658, N1505);
nor NOR2 (N2674, N2667, N2129);
and AND2 (N2675, N2673, N2136);
not NOT1 (N2676, N2670);
nand NAND3 (N2677, N2671, N2596, N1547);
nor NOR4 (N2678, N2677, N254, N1417, N1976);
nand NAND2 (N2679, N2672, N1349);
nor NOR3 (N2680, N2674, N1917, N2637);
nand NAND3 (N2681, N2669, N793, N604);
or OR2 (N2682, N2662, N476);
not NOT1 (N2683, N2675);
not NOT1 (N2684, N2678);
or OR4 (N2685, N2679, N1242, N2586, N1556);
buf BUF1 (N2686, N2685);
nand NAND4 (N2687, N2686, N2403, N1536, N1683);
xor XOR2 (N2688, N2684, N1680);
not NOT1 (N2689, N2625);
xor XOR2 (N2690, N2680, N256);
buf BUF1 (N2691, N2688);
nor NOR4 (N2692, N2666, N654, N1212, N2526);
and AND2 (N2693, N2689, N485);
or OR2 (N2694, N2682, N1448);
not NOT1 (N2695, N2681);
nand NAND4 (N2696, N2691, N903, N1728, N2108);
and AND4 (N2697, N2692, N735, N1541, N1090);
not NOT1 (N2698, N2668);
or OR4 (N2699, N2697, N263, N2120, N315);
not NOT1 (N2700, N2693);
xor XOR2 (N2701, N2699, N2256);
buf BUF1 (N2702, N2676);
or OR4 (N2703, N2683, N284, N1537, N2);
nor NOR3 (N2704, N2700, N1231, N1535);
nand NAND2 (N2705, N2701, N769);
and AND4 (N2706, N2703, N642, N2549, N694);
buf BUF1 (N2707, N2702);
not NOT1 (N2708, N2690);
and AND3 (N2709, N2698, N376, N1930);
xor XOR2 (N2710, N2705, N920);
and AND4 (N2711, N2696, N2689, N2321, N797);
buf BUF1 (N2712, N2695);
nor NOR4 (N2713, N2706, N107, N287, N1778);
buf BUF1 (N2714, N2712);
or OR4 (N2715, N2704, N2189, N841, N2507);
and AND3 (N2716, N2709, N329, N570);
not NOT1 (N2717, N2711);
xor XOR2 (N2718, N2710, N128);
xor XOR2 (N2719, N2716, N1110);
xor XOR2 (N2720, N2687, N2567);
or OR4 (N2721, N2708, N759, N1716, N2080);
nand NAND2 (N2722, N2715, N331);
not NOT1 (N2723, N2714);
not NOT1 (N2724, N2694);
and AND3 (N2725, N2718, N984, N559);
not NOT1 (N2726, N2717);
not NOT1 (N2727, N2713);
buf BUF1 (N2728, N2725);
xor XOR2 (N2729, N2728, N520);
not NOT1 (N2730, N2719);
buf BUF1 (N2731, N2726);
buf BUF1 (N2732, N2729);
not NOT1 (N2733, N2731);
or OR2 (N2734, N2732, N1729);
nor NOR4 (N2735, N2723, N1623, N1466, N1545);
nor NOR3 (N2736, N2722, N2288, N367);
or OR2 (N2737, N2733, N1832);
not NOT1 (N2738, N2734);
and AND4 (N2739, N2735, N2081, N926, N1037);
nand NAND4 (N2740, N2724, N1777, N2158, N717);
xor XOR2 (N2741, N2727, N2124);
xor XOR2 (N2742, N2740, N2208);
buf BUF1 (N2743, N2707);
not NOT1 (N2744, N2737);
not NOT1 (N2745, N2742);
and AND4 (N2746, N2721, N2421, N838, N399);
buf BUF1 (N2747, N2730);
or OR2 (N2748, N2738, N797);
xor XOR2 (N2749, N2743, N407);
buf BUF1 (N2750, N2744);
or OR2 (N2751, N2739, N511);
nor NOR3 (N2752, N2749, N48, N1816);
nor NOR2 (N2753, N2752, N1497);
buf BUF1 (N2754, N2750);
not NOT1 (N2755, N2748);
not NOT1 (N2756, N2751);
not NOT1 (N2757, N2756);
nand NAND2 (N2758, N2736, N1545);
xor XOR2 (N2759, N2746, N494);
not NOT1 (N2760, N2754);
xor XOR2 (N2761, N2760, N546);
nand NAND3 (N2762, N2745, N890, N1597);
not NOT1 (N2763, N2755);
or OR3 (N2764, N2741, N1046, N1592);
or OR2 (N2765, N2761, N480);
and AND3 (N2766, N2762, N382, N2722);
nand NAND4 (N2767, N2765, N1478, N230, N1511);
not NOT1 (N2768, N2764);
nand NAND4 (N2769, N2758, N1240, N1810, N1999);
or OR4 (N2770, N2763, N2065, N1859, N2495);
nand NAND2 (N2771, N2720, N1256);
and AND3 (N2772, N2747, N610, N294);
nand NAND2 (N2773, N2757, N1615);
nor NOR4 (N2774, N2767, N863, N721, N1185);
and AND3 (N2775, N2769, N2006, N231);
buf BUF1 (N2776, N2766);
not NOT1 (N2777, N2775);
buf BUF1 (N2778, N2774);
and AND2 (N2779, N2771, N820);
or OR4 (N2780, N2770, N449, N2703, N698);
not NOT1 (N2781, N2753);
nor NOR4 (N2782, N2776, N1412, N76, N2196);
buf BUF1 (N2783, N2782);
or OR4 (N2784, N2780, N1786, N2068, N2742);
or OR3 (N2785, N2759, N1711, N464);
not NOT1 (N2786, N2773);
xor XOR2 (N2787, N2786, N950);
xor XOR2 (N2788, N2778, N2235);
xor XOR2 (N2789, N2783, N860);
and AND4 (N2790, N2785, N2575, N589, N1195);
nor NOR4 (N2791, N2784, N1945, N1182, N719);
and AND2 (N2792, N2777, N813);
nor NOR3 (N2793, N2787, N1895, N1324);
and AND3 (N2794, N2790, N1198, N437);
and AND2 (N2795, N2793, N1111);
not NOT1 (N2796, N2768);
and AND3 (N2797, N2789, N1799, N822);
not NOT1 (N2798, N2792);
xor XOR2 (N2799, N2779, N557);
nand NAND2 (N2800, N2781, N1421);
and AND2 (N2801, N2772, N2148);
or OR4 (N2802, N2799, N2700, N1044, N1969);
or OR4 (N2803, N2796, N2268, N230, N2739);
or OR2 (N2804, N2791, N1326);
nand NAND4 (N2805, N2794, N2797, N445, N70);
and AND4 (N2806, N286, N1457, N185, N1089);
nor NOR3 (N2807, N2806, N459, N946);
nand NAND3 (N2808, N2803, N1512, N2394);
or OR4 (N2809, N2808, N1361, N1727, N739);
buf BUF1 (N2810, N2801);
buf BUF1 (N2811, N2807);
buf BUF1 (N2812, N2811);
buf BUF1 (N2813, N2812);
nand NAND3 (N2814, N2805, N989, N2217);
or OR3 (N2815, N2795, N808, N473);
buf BUF1 (N2816, N2804);
and AND4 (N2817, N2788, N573, N1475, N1853);
and AND4 (N2818, N2815, N758, N1653, N349);
nor NOR2 (N2819, N2817, N2294);
nor NOR3 (N2820, N2816, N2794, N1597);
nand NAND2 (N2821, N2798, N1756);
not NOT1 (N2822, N2814);
xor XOR2 (N2823, N2820, N1193);
nor NOR3 (N2824, N2823, N27, N2756);
and AND3 (N2825, N2822, N2719, N58);
nor NOR4 (N2826, N2810, N2466, N2371, N1801);
and AND3 (N2827, N2819, N492, N1097);
buf BUF1 (N2828, N2826);
not NOT1 (N2829, N2802);
xor XOR2 (N2830, N2821, N86);
nor NOR4 (N2831, N2829, N108, N18, N1135);
or OR4 (N2832, N2830, N1117, N892, N1248);
not NOT1 (N2833, N2809);
buf BUF1 (N2834, N2832);
buf BUF1 (N2835, N2833);
or OR3 (N2836, N2818, N1017, N2136);
or OR3 (N2837, N2827, N2103, N709);
not NOT1 (N2838, N2834);
nor NOR3 (N2839, N2838, N1663, N1454);
not NOT1 (N2840, N2828);
and AND4 (N2841, N2825, N2513, N2027, N317);
xor XOR2 (N2842, N2841, N2024);
nand NAND2 (N2843, N2840, N2153);
or OR3 (N2844, N2839, N1620, N1995);
and AND4 (N2845, N2813, N1698, N1532, N2263);
not NOT1 (N2846, N2842);
xor XOR2 (N2847, N2845, N225);
buf BUF1 (N2848, N2846);
or OR2 (N2849, N2837, N2582);
xor XOR2 (N2850, N2800, N2177);
nand NAND3 (N2851, N2848, N237, N1162);
and AND2 (N2852, N2824, N213);
or OR2 (N2853, N2847, N1698);
and AND3 (N2854, N2836, N2070, N237);
or OR4 (N2855, N2851, N131, N1838, N396);
or OR2 (N2856, N2852, N1048);
xor XOR2 (N2857, N2855, N42);
xor XOR2 (N2858, N2831, N651);
and AND3 (N2859, N2853, N1074, N2603);
buf BUF1 (N2860, N2856);
nor NOR4 (N2861, N2850, N527, N2507, N1257);
xor XOR2 (N2862, N2849, N2142);
nor NOR3 (N2863, N2854, N2324, N712);
xor XOR2 (N2864, N2862, N1321);
nand NAND4 (N2865, N2863, N1291, N2583, N1788);
and AND3 (N2866, N2860, N1032, N1364);
or OR4 (N2867, N2858, N1806, N948, N2155);
or OR4 (N2868, N2861, N1887, N2004, N2414);
buf BUF1 (N2869, N2857);
and AND3 (N2870, N2868, N2227, N826);
or OR3 (N2871, N2859, N1422, N2368);
nand NAND2 (N2872, N2865, N598);
buf BUF1 (N2873, N2869);
nor NOR4 (N2874, N2871, N2767, N1170, N1063);
not NOT1 (N2875, N2870);
not NOT1 (N2876, N2867);
xor XOR2 (N2877, N2835, N1075);
and AND4 (N2878, N2864, N1197, N1670, N2610);
and AND3 (N2879, N2878, N1255, N1041);
and AND4 (N2880, N2876, N2660, N592, N1361);
nand NAND2 (N2881, N2874, N2521);
buf BUF1 (N2882, N2880);
and AND2 (N2883, N2879, N239);
buf BUF1 (N2884, N2844);
not NOT1 (N2885, N2884);
xor XOR2 (N2886, N2881, N432);
or OR2 (N2887, N2883, N1100);
or OR4 (N2888, N2877, N1422, N305, N2423);
or OR2 (N2889, N2873, N724);
or OR4 (N2890, N2875, N2139, N1834, N325);
xor XOR2 (N2891, N2888, N2402);
and AND2 (N2892, N2891, N1668);
buf BUF1 (N2893, N2892);
nand NAND3 (N2894, N2886, N2691, N440);
or OR4 (N2895, N2843, N463, N1835, N725);
or OR4 (N2896, N2895, N7, N2339, N2668);
and AND2 (N2897, N2882, N2654);
xor XOR2 (N2898, N2896, N2417);
and AND3 (N2899, N2872, N2714, N920);
xor XOR2 (N2900, N2898, N2418);
and AND3 (N2901, N2866, N913, N764);
and AND4 (N2902, N2901, N333, N89, N1668);
or OR2 (N2903, N2899, N2629);
nor NOR3 (N2904, N2889, N1672, N2346);
not NOT1 (N2905, N2902);
and AND3 (N2906, N2890, N1937, N1668);
xor XOR2 (N2907, N2903, N2536);
xor XOR2 (N2908, N2897, N1369);
nand NAND2 (N2909, N2893, N2692);
buf BUF1 (N2910, N2900);
or OR4 (N2911, N2885, N1197, N638, N2705);
nor NOR3 (N2912, N2909, N256, N2509);
nor NOR4 (N2913, N2910, N2760, N1900, N1922);
nor NOR4 (N2914, N2913, N2096, N686, N962);
or OR3 (N2915, N2911, N1877, N642);
nor NOR3 (N2916, N2907, N2743, N236);
buf BUF1 (N2917, N2915);
or OR2 (N2918, N2904, N69);
not NOT1 (N2919, N2894);
nor NOR4 (N2920, N2912, N429, N2110, N1020);
nand NAND2 (N2921, N2905, N1303);
or OR3 (N2922, N2920, N442, N2237);
buf BUF1 (N2923, N2887);
and AND2 (N2924, N2906, N206);
buf BUF1 (N2925, N2918);
xor XOR2 (N2926, N2924, N2073);
not NOT1 (N2927, N2919);
and AND4 (N2928, N2908, N2728, N2832, N2448);
xor XOR2 (N2929, N2917, N1885);
buf BUF1 (N2930, N2926);
and AND2 (N2931, N2925, N1009);
xor XOR2 (N2932, N2922, N1777);
nand NAND2 (N2933, N2931, N1445);
nand NAND4 (N2934, N2933, N2655, N366, N2166);
nor NOR3 (N2935, N2921, N2367, N1862);
nor NOR3 (N2936, N2916, N1783, N630);
or OR3 (N2937, N2929, N136, N1820);
not NOT1 (N2938, N2927);
buf BUF1 (N2939, N2932);
buf BUF1 (N2940, N2914);
and AND4 (N2941, N2935, N1239, N1336, N2425);
and AND2 (N2942, N2940, N383);
and AND2 (N2943, N2938, N2862);
nand NAND3 (N2944, N2937, N1706, N2674);
and AND3 (N2945, N2941, N1225, N1563);
buf BUF1 (N2946, N2923);
nor NOR2 (N2947, N2936, N554);
and AND2 (N2948, N2947, N842);
and AND4 (N2949, N2942, N151, N1679, N9);
nor NOR2 (N2950, N2949, N1061);
xor XOR2 (N2951, N2944, N482);
and AND3 (N2952, N2950, N414, N349);
buf BUF1 (N2953, N2945);
and AND4 (N2954, N2948, N791, N1058, N2781);
nor NOR2 (N2955, N2934, N1580);
and AND2 (N2956, N2930, N1239);
nand NAND2 (N2957, N2928, N815);
nor NOR4 (N2958, N2953, N1015, N1267, N1160);
buf BUF1 (N2959, N2943);
or OR3 (N2960, N2957, N181, N2718);
or OR4 (N2961, N2956, N2155, N1936, N2623);
not NOT1 (N2962, N2954);
nor NOR3 (N2963, N2962, N107, N343);
not NOT1 (N2964, N2961);
nor NOR4 (N2965, N2946, N166, N568, N2536);
and AND3 (N2966, N2955, N1482, N1763);
or OR2 (N2967, N2964, N1374);
or OR3 (N2968, N2967, N2037, N1758);
xor XOR2 (N2969, N2966, N2284);
not NOT1 (N2970, N2958);
or OR4 (N2971, N2968, N2785, N1194, N1115);
not NOT1 (N2972, N2960);
nand NAND4 (N2973, N2970, N2301, N1470, N1635);
and AND3 (N2974, N2971, N502, N2839);
xor XOR2 (N2975, N2969, N1266);
nand NAND3 (N2976, N2939, N2578, N939);
xor XOR2 (N2977, N2963, N1591);
not NOT1 (N2978, N2974);
not NOT1 (N2979, N2951);
nand NAND2 (N2980, N2965, N1086);
or OR3 (N2981, N2972, N1272, N1964);
buf BUF1 (N2982, N2977);
nor NOR2 (N2983, N2980, N716);
nand NAND3 (N2984, N2982, N1841, N1731);
and AND3 (N2985, N2979, N1914, N2574);
nand NAND2 (N2986, N2985, N1257);
buf BUF1 (N2987, N2975);
nand NAND2 (N2988, N2976, N927);
nand NAND3 (N2989, N2952, N2095, N1060);
buf BUF1 (N2990, N2989);
and AND3 (N2991, N2978, N2380, N565);
xor XOR2 (N2992, N2988, N2920);
nand NAND2 (N2993, N2984, N15);
and AND3 (N2994, N2993, N2278, N1544);
or OR3 (N2995, N2986, N2867, N2444);
nand NAND2 (N2996, N2981, N961);
xor XOR2 (N2997, N2992, N358);
and AND3 (N2998, N2994, N2195, N883);
nor NOR2 (N2999, N2998, N383);
nand NAND3 (N3000, N2995, N1537, N2604);
or OR3 (N3001, N2991, N1180, N855);
xor XOR2 (N3002, N2987, N391);
nor NOR2 (N3003, N2999, N1348);
nand NAND4 (N3004, N2959, N2348, N987, N976);
or OR4 (N3005, N3004, N2329, N253, N1754);
xor XOR2 (N3006, N3001, N2317);
not NOT1 (N3007, N2990);
or OR3 (N3008, N2973, N2189, N2815);
nor NOR3 (N3009, N2997, N1289, N929);
xor XOR2 (N3010, N3002, N1936);
buf BUF1 (N3011, N3009);
buf BUF1 (N3012, N3000);
buf BUF1 (N3013, N3007);
endmodule