// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10;

output N608,N596,N606,N609,N605,N607,N587,N594,N597,N610;

and AND4 (N11, N8, N3, N5, N6);
nor NOR4 (N12, N1, N3, N7, N9);
and AND3 (N13, N2, N12, N12);
or OR3 (N14, N10, N2, N12);
nor NOR3 (N15, N3, N4, N11);
xor XOR2 (N16, N14, N5);
buf BUF1 (N17, N5);
not NOT1 (N18, N4);
xor XOR2 (N19, N8, N15);
nand NAND2 (N20, N3, N6);
buf BUF1 (N21, N17);
and AND4 (N22, N7, N6, N5, N12);
or OR2 (N23, N10, N20);
not NOT1 (N24, N2);
xor XOR2 (N25, N20, N20);
xor XOR2 (N26, N7, N18);
and AND2 (N27, N22, N22);
nand NAND2 (N28, N15, N23);
not NOT1 (N29, N27);
nand NAND2 (N30, N13, N5);
nor NOR4 (N31, N26, N5, N17, N18);
buf BUF1 (N32, N2);
or OR4 (N33, N30, N10, N11, N8);
xor XOR2 (N34, N21, N12);
nand NAND2 (N35, N16, N33);
nor NOR4 (N36, N14, N32, N21, N25);
nand NAND3 (N37, N7, N23, N1);
or OR4 (N38, N17, N7, N33, N6);
nand NAND3 (N39, N31, N3, N25);
not NOT1 (N40, N38);
and AND2 (N41, N37, N11);
nand NAND2 (N42, N28, N12);
not NOT1 (N43, N39);
not NOT1 (N44, N19);
and AND2 (N45, N24, N27);
not NOT1 (N46, N40);
and AND4 (N47, N35, N10, N16, N21);
not NOT1 (N48, N36);
not NOT1 (N49, N44);
nand NAND2 (N50, N41, N47);
buf BUF1 (N51, N50);
xor XOR2 (N52, N23, N18);
buf BUF1 (N53, N52);
and AND4 (N54, N49, N49, N29, N10);
nand NAND3 (N55, N34, N53, N17);
nand NAND2 (N56, N29, N54);
nor NOR2 (N57, N10, N34);
or OR2 (N58, N16, N10);
or OR2 (N59, N45, N25);
nor NOR4 (N60, N59, N45, N7, N18);
nor NOR3 (N61, N56, N55, N33);
not NOT1 (N62, N32);
or OR3 (N63, N60, N59, N2);
not NOT1 (N64, N62);
and AND3 (N65, N51, N52, N23);
buf BUF1 (N66, N58);
buf BUF1 (N67, N57);
and AND3 (N68, N67, N16, N1);
buf BUF1 (N69, N64);
and AND4 (N70, N68, N32, N45, N26);
nand NAND3 (N71, N70, N45, N39);
and AND2 (N72, N65, N22);
buf BUF1 (N73, N43);
nor NOR2 (N74, N63, N57);
buf BUF1 (N75, N71);
buf BUF1 (N76, N69);
and AND4 (N77, N42, N15, N26, N37);
xor XOR2 (N78, N77, N22);
or OR4 (N79, N61, N41, N21, N4);
xor XOR2 (N80, N66, N7);
not NOT1 (N81, N78);
and AND4 (N82, N81, N77, N53, N33);
nand NAND3 (N83, N82, N52, N15);
nor NOR4 (N84, N79, N60, N15, N34);
buf BUF1 (N85, N48);
nand NAND2 (N86, N73, N64);
not NOT1 (N87, N46);
nor NOR4 (N88, N87, N64, N39, N59);
nor NOR3 (N89, N76, N22, N83);
buf BUF1 (N90, N37);
or OR3 (N91, N90, N64, N65);
not NOT1 (N92, N74);
not NOT1 (N93, N92);
not NOT1 (N94, N80);
not NOT1 (N95, N84);
buf BUF1 (N96, N94);
buf BUF1 (N97, N75);
nand NAND4 (N98, N95, N70, N52, N63);
nor NOR4 (N99, N85, N39, N98, N20);
nand NAND2 (N100, N96, N30);
not NOT1 (N101, N62);
not NOT1 (N102, N86);
nor NOR3 (N103, N97, N2, N101);
nand NAND4 (N104, N20, N33, N85, N16);
xor XOR2 (N105, N104, N61);
not NOT1 (N106, N103);
xor XOR2 (N107, N88, N19);
and AND2 (N108, N89, N28);
buf BUF1 (N109, N72);
and AND3 (N110, N99, N11, N72);
nand NAND4 (N111, N93, N38, N106, N33);
xor XOR2 (N112, N8, N16);
not NOT1 (N113, N105);
not NOT1 (N114, N113);
and AND2 (N115, N100, N27);
buf BUF1 (N116, N112);
xor XOR2 (N117, N109, N30);
and AND2 (N118, N91, N2);
or OR2 (N119, N108, N110);
nand NAND4 (N120, N55, N31, N98, N83);
not NOT1 (N121, N117);
buf BUF1 (N122, N120);
not NOT1 (N123, N119);
nand NAND4 (N124, N102, N101, N117, N102);
xor XOR2 (N125, N107, N29);
xor XOR2 (N126, N121, N118);
and AND3 (N127, N11, N19, N120);
or OR2 (N128, N122, N3);
xor XOR2 (N129, N115, N124);
nand NAND3 (N130, N108, N118, N35);
and AND3 (N131, N129, N112, N11);
xor XOR2 (N132, N126, N6);
nor NOR4 (N133, N132, N43, N83, N81);
not NOT1 (N134, N131);
nand NAND4 (N135, N133, N100, N66, N126);
xor XOR2 (N136, N114, N95);
not NOT1 (N137, N136);
buf BUF1 (N138, N135);
buf BUF1 (N139, N138);
xor XOR2 (N140, N128, N32);
and AND4 (N141, N123, N138, N113, N11);
nand NAND4 (N142, N127, N66, N88, N22);
nand NAND3 (N143, N137, N68, N97);
or OR2 (N144, N134, N132);
nor NOR2 (N145, N139, N34);
buf BUF1 (N146, N130);
or OR3 (N147, N111, N86, N30);
not NOT1 (N148, N144);
not NOT1 (N149, N147);
xor XOR2 (N150, N140, N113);
not NOT1 (N151, N143);
or OR4 (N152, N149, N91, N48, N95);
nor NOR3 (N153, N152, N138, N21);
nor NOR2 (N154, N146, N134);
not NOT1 (N155, N148);
xor XOR2 (N156, N154, N79);
nand NAND3 (N157, N116, N43, N135);
and AND3 (N158, N150, N6, N136);
xor XOR2 (N159, N141, N149);
nor NOR2 (N160, N158, N7);
not NOT1 (N161, N142);
and AND2 (N162, N151, N24);
or OR4 (N163, N156, N160, N5, N47);
xor XOR2 (N164, N105, N24);
xor XOR2 (N165, N125, N134);
and AND3 (N166, N145, N93, N58);
nand NAND2 (N167, N165, N105);
and AND2 (N168, N157, N99);
nor NOR3 (N169, N163, N15, N121);
xor XOR2 (N170, N164, N148);
nor NOR2 (N171, N170, N22);
or OR3 (N172, N159, N119, N46);
nand NAND4 (N173, N168, N7, N27, N113);
buf BUF1 (N174, N167);
xor XOR2 (N175, N171, N120);
nand NAND4 (N176, N153, N113, N75, N75);
nand NAND2 (N177, N161, N113);
or OR2 (N178, N155, N19);
or OR2 (N179, N166, N96);
and AND4 (N180, N174, N130, N106, N165);
and AND2 (N181, N175, N1);
nor NOR2 (N182, N162, N31);
or OR2 (N183, N173, N46);
nor NOR4 (N184, N182, N150, N22, N179);
xor XOR2 (N185, N157, N115);
not NOT1 (N186, N177);
nand NAND4 (N187, N183, N1, N115, N51);
nand NAND2 (N188, N172, N47);
not NOT1 (N189, N186);
xor XOR2 (N190, N169, N188);
xor XOR2 (N191, N112, N78);
buf BUF1 (N192, N178);
nand NAND2 (N193, N191, N129);
nand NAND2 (N194, N189, N187);
not NOT1 (N195, N38);
xor XOR2 (N196, N192, N146);
or OR2 (N197, N176, N169);
buf BUF1 (N198, N185);
or OR3 (N199, N193, N59, N20);
not NOT1 (N200, N194);
nand NAND4 (N201, N190, N156, N52, N128);
buf BUF1 (N202, N181);
xor XOR2 (N203, N184, N158);
buf BUF1 (N204, N200);
nand NAND2 (N205, N203, N39);
or OR4 (N206, N205, N127, N119, N114);
buf BUF1 (N207, N197);
buf BUF1 (N208, N180);
not NOT1 (N209, N198);
and AND4 (N210, N196, N147, N11, N44);
and AND3 (N211, N202, N197, N96);
xor XOR2 (N212, N206, N116);
not NOT1 (N213, N209);
buf BUF1 (N214, N212);
or OR2 (N215, N204, N59);
buf BUF1 (N216, N215);
nor NOR4 (N217, N195, N115, N199, N201);
not NOT1 (N218, N139);
xor XOR2 (N219, N167, N123);
not NOT1 (N220, N210);
and AND2 (N221, N214, N72);
and AND3 (N222, N216, N179, N181);
buf BUF1 (N223, N219);
nand NAND4 (N224, N213, N52, N117, N141);
xor XOR2 (N225, N217, N168);
or OR2 (N226, N218, N143);
buf BUF1 (N227, N220);
xor XOR2 (N228, N211, N115);
buf BUF1 (N229, N208);
not NOT1 (N230, N223);
nor NOR3 (N231, N227, N112, N223);
nor NOR2 (N232, N225, N112);
not NOT1 (N233, N224);
nor NOR3 (N234, N233, N16, N119);
buf BUF1 (N235, N234);
or OR3 (N236, N207, N80, N81);
buf BUF1 (N237, N226);
not NOT1 (N238, N237);
or OR3 (N239, N228, N43, N150);
nand NAND3 (N240, N229, N57, N79);
not NOT1 (N241, N222);
nor NOR4 (N242, N231, N48, N38, N229);
and AND3 (N243, N239, N224, N224);
nor NOR3 (N244, N236, N208, N15);
xor XOR2 (N245, N232, N216);
xor XOR2 (N246, N238, N174);
nand NAND3 (N247, N242, N29, N69);
nand NAND2 (N248, N247, N188);
nand NAND4 (N249, N245, N71, N36, N201);
nor NOR4 (N250, N248, N224, N230, N65);
not NOT1 (N251, N134);
buf BUF1 (N252, N246);
xor XOR2 (N253, N243, N190);
or OR2 (N254, N251, N107);
not NOT1 (N255, N240);
nand NAND3 (N256, N254, N225, N29);
xor XOR2 (N257, N256, N38);
not NOT1 (N258, N241);
and AND4 (N259, N249, N173, N128, N44);
and AND4 (N260, N253, N194, N100, N17);
xor XOR2 (N261, N257, N125);
nand NAND3 (N262, N221, N35, N47);
or OR3 (N263, N235, N42, N166);
or OR3 (N264, N252, N261, N93);
nor NOR4 (N265, N223, N44, N262, N11);
not NOT1 (N266, N18);
xor XOR2 (N267, N264, N254);
or OR3 (N268, N267, N35, N137);
and AND4 (N269, N258, N238, N63, N126);
buf BUF1 (N270, N250);
nor NOR3 (N271, N265, N244, N136);
not NOT1 (N272, N18);
nand NAND2 (N273, N268, N153);
not NOT1 (N274, N273);
and AND3 (N275, N270, N244, N254);
not NOT1 (N276, N255);
and AND2 (N277, N266, N216);
and AND4 (N278, N271, N201, N209, N201);
and AND2 (N279, N259, N120);
or OR2 (N280, N279, N140);
buf BUF1 (N281, N263);
or OR4 (N282, N260, N229, N6, N231);
not NOT1 (N283, N276);
and AND2 (N284, N280, N271);
buf BUF1 (N285, N269);
and AND3 (N286, N282, N209, N52);
buf BUF1 (N287, N278);
nor NOR2 (N288, N272, N52);
xor XOR2 (N289, N274, N204);
buf BUF1 (N290, N284);
xor XOR2 (N291, N287, N87);
buf BUF1 (N292, N286);
nor NOR4 (N293, N275, N141, N119, N69);
buf BUF1 (N294, N291);
xor XOR2 (N295, N277, N199);
and AND2 (N296, N289, N30);
nor NOR2 (N297, N292, N48);
buf BUF1 (N298, N295);
nand NAND2 (N299, N296, N196);
and AND3 (N300, N294, N131, N246);
and AND2 (N301, N285, N167);
nand NAND2 (N302, N281, N237);
nand NAND2 (N303, N299, N215);
nor NOR3 (N304, N297, N33, N259);
nand NAND2 (N305, N301, N187);
xor XOR2 (N306, N303, N26);
nor NOR2 (N307, N306, N265);
nand NAND2 (N308, N307, N201);
xor XOR2 (N309, N308, N288);
or OR3 (N310, N290, N304, N176);
xor XOR2 (N311, N118, N43);
buf BUF1 (N312, N147);
xor XOR2 (N313, N293, N209);
xor XOR2 (N314, N312, N65);
not NOT1 (N315, N314);
nand NAND2 (N316, N310, N109);
nand NAND3 (N317, N311, N111, N149);
buf BUF1 (N318, N298);
nor NOR3 (N319, N302, N16, N188);
buf BUF1 (N320, N319);
buf BUF1 (N321, N320);
and AND3 (N322, N305, N133, N55);
xor XOR2 (N323, N322, N45);
nor NOR3 (N324, N300, N157, N309);
and AND4 (N325, N6, N217, N229, N105);
xor XOR2 (N326, N316, N98);
and AND2 (N327, N315, N201);
nor NOR3 (N328, N324, N146, N257);
nand NAND3 (N329, N318, N199, N143);
xor XOR2 (N330, N327, N268);
not NOT1 (N331, N283);
xor XOR2 (N332, N328, N152);
nand NAND4 (N333, N323, N285, N209, N265);
buf BUF1 (N334, N331);
nor NOR4 (N335, N330, N31, N199, N283);
not NOT1 (N336, N325);
not NOT1 (N337, N335);
xor XOR2 (N338, N336, N261);
nand NAND2 (N339, N317, N316);
buf BUF1 (N340, N332);
not NOT1 (N341, N340);
and AND2 (N342, N337, N270);
or OR3 (N343, N334, N52, N147);
and AND4 (N344, N341, N330, N311, N13);
not NOT1 (N345, N343);
not NOT1 (N346, N339);
not NOT1 (N347, N338);
buf BUF1 (N348, N329);
buf BUF1 (N349, N313);
nor NOR3 (N350, N347, N199, N263);
and AND4 (N351, N321, N8, N126, N340);
and AND4 (N352, N345, N25, N7, N253);
and AND4 (N353, N352, N9, N247, N224);
nand NAND2 (N354, N342, N75);
xor XOR2 (N355, N351, N235);
buf BUF1 (N356, N348);
and AND2 (N357, N344, N99);
buf BUF1 (N358, N357);
buf BUF1 (N359, N326);
and AND2 (N360, N354, N251);
nor NOR2 (N361, N353, N203);
xor XOR2 (N362, N355, N239);
nand NAND3 (N363, N360, N153, N20);
buf BUF1 (N364, N333);
xor XOR2 (N365, N350, N326);
and AND4 (N366, N362, N360, N195, N57);
and AND2 (N367, N358, N169);
nor NOR3 (N368, N364, N62, N53);
xor XOR2 (N369, N359, N239);
xor XOR2 (N370, N368, N323);
xor XOR2 (N371, N356, N246);
nor NOR4 (N372, N371, N51, N53, N303);
nor NOR4 (N373, N372, N249, N80, N161);
xor XOR2 (N374, N366, N10);
and AND2 (N375, N346, N148);
or OR3 (N376, N365, N161, N8);
buf BUF1 (N377, N374);
and AND2 (N378, N377, N349);
or OR3 (N379, N378, N129, N93);
xor XOR2 (N380, N286, N102);
xor XOR2 (N381, N363, N61);
nor NOR3 (N382, N373, N227, N240);
nor NOR3 (N383, N380, N100, N180);
xor XOR2 (N384, N382, N321);
nand NAND2 (N385, N369, N65);
nor NOR2 (N386, N384, N42);
not NOT1 (N387, N367);
buf BUF1 (N388, N385);
or OR3 (N389, N376, N233, N220);
nor NOR3 (N390, N381, N159, N36);
nor NOR3 (N391, N389, N31, N256);
and AND4 (N392, N390, N14, N247, N89);
or OR4 (N393, N386, N37, N141, N33);
buf BUF1 (N394, N393);
not NOT1 (N395, N387);
buf BUF1 (N396, N375);
buf BUF1 (N397, N391);
and AND4 (N398, N397, N146, N134, N207);
nand NAND3 (N399, N392, N55, N11);
and AND2 (N400, N398, N93);
not NOT1 (N401, N388);
not NOT1 (N402, N370);
not NOT1 (N403, N383);
nand NAND4 (N404, N399, N165, N194, N335);
and AND3 (N405, N361, N201, N77);
not NOT1 (N406, N394);
nor NOR3 (N407, N396, N42, N25);
and AND4 (N408, N403, N329, N165, N89);
nor NOR4 (N409, N401, N14, N98, N3);
or OR2 (N410, N405, N354);
nand NAND4 (N411, N406, N404, N9, N327);
not NOT1 (N412, N176);
xor XOR2 (N413, N411, N169);
or OR2 (N414, N413, N344);
nor NOR2 (N415, N408, N179);
buf BUF1 (N416, N414);
nand NAND4 (N417, N407, N314, N51, N15);
or OR3 (N418, N395, N243, N333);
buf BUF1 (N419, N416);
or OR3 (N420, N409, N307, N325);
buf BUF1 (N421, N420);
and AND4 (N422, N412, N92, N117, N32);
or OR4 (N423, N402, N338, N325, N288);
buf BUF1 (N424, N379);
xor XOR2 (N425, N421, N84);
not NOT1 (N426, N410);
and AND2 (N427, N417, N124);
buf BUF1 (N428, N400);
or OR4 (N429, N418, N238, N263, N109);
not NOT1 (N430, N423);
nand NAND2 (N431, N426, N300);
not NOT1 (N432, N424);
nor NOR2 (N433, N419, N411);
not NOT1 (N434, N430);
nor NOR4 (N435, N422, N56, N420, N254);
xor XOR2 (N436, N434, N256);
nand NAND2 (N437, N436, N240);
nor NOR3 (N438, N433, N143, N428);
buf BUF1 (N439, N340);
buf BUF1 (N440, N425);
or OR2 (N441, N438, N361);
or OR4 (N442, N432, N353, N262, N1);
not NOT1 (N443, N435);
buf BUF1 (N444, N431);
and AND3 (N445, N427, N306, N50);
xor XOR2 (N446, N415, N355);
and AND3 (N447, N441, N443, N30);
xor XOR2 (N448, N388, N400);
and AND2 (N449, N437, N91);
not NOT1 (N450, N446);
buf BUF1 (N451, N444);
nand NAND4 (N452, N450, N28, N303, N23);
and AND2 (N453, N439, N78);
and AND2 (N454, N452, N371);
not NOT1 (N455, N429);
nand NAND2 (N456, N442, N129);
nor NOR2 (N457, N453, N271);
nor NOR2 (N458, N455, N328);
nor NOR3 (N459, N451, N86, N448);
not NOT1 (N460, N16);
buf BUF1 (N461, N454);
nand NAND3 (N462, N456, N46, N75);
buf BUF1 (N463, N445);
and AND4 (N464, N449, N247, N54, N395);
nor NOR3 (N465, N459, N108, N239);
not NOT1 (N466, N458);
xor XOR2 (N467, N466, N36);
xor XOR2 (N468, N464, N330);
and AND2 (N469, N440, N262);
not NOT1 (N470, N457);
xor XOR2 (N471, N447, N371);
not NOT1 (N472, N465);
and AND3 (N473, N472, N22, N317);
buf BUF1 (N474, N470);
or OR2 (N475, N474, N330);
buf BUF1 (N476, N471);
nand NAND4 (N477, N468, N213, N310, N251);
and AND2 (N478, N473, N298);
or OR4 (N479, N467, N355, N432, N114);
xor XOR2 (N480, N463, N74);
and AND4 (N481, N476, N246, N354, N134);
and AND4 (N482, N479, N396, N109, N348);
xor XOR2 (N483, N469, N214);
and AND2 (N484, N481, N399);
nor NOR2 (N485, N461, N77);
nor NOR3 (N486, N478, N376, N73);
not NOT1 (N487, N477);
or OR4 (N488, N486, N485, N399, N191);
not NOT1 (N489, N108);
nor NOR4 (N490, N475, N137, N269, N363);
or OR4 (N491, N482, N86, N106, N170);
or OR3 (N492, N489, N258, N360);
xor XOR2 (N493, N487, N115);
or OR2 (N494, N480, N67);
nor NOR2 (N495, N462, N383);
nand NAND2 (N496, N492, N446);
nand NAND4 (N497, N488, N210, N460, N458);
nor NOR4 (N498, N246, N67, N342, N342);
or OR3 (N499, N491, N297, N378);
or OR3 (N500, N498, N271, N230);
nand NAND3 (N501, N499, N458, N68);
not NOT1 (N502, N484);
nor NOR2 (N503, N497, N162);
and AND2 (N504, N501, N46);
or OR3 (N505, N496, N305, N163);
xor XOR2 (N506, N494, N56);
or OR4 (N507, N502, N158, N177, N84);
or OR3 (N508, N490, N6, N16);
or OR3 (N509, N505, N37, N146);
or OR2 (N510, N507, N319);
or OR4 (N511, N506, N195, N372, N222);
or OR2 (N512, N483, N212);
nand NAND2 (N513, N509, N497);
buf BUF1 (N514, N513);
xor XOR2 (N515, N504, N361);
or OR2 (N516, N514, N428);
nor NOR2 (N517, N516, N236);
or OR4 (N518, N500, N202, N31, N236);
nand NAND2 (N519, N508, N461);
and AND4 (N520, N517, N16, N186, N439);
and AND3 (N521, N510, N352, N380);
nor NOR2 (N522, N520, N455);
xor XOR2 (N523, N511, N411);
xor XOR2 (N524, N512, N143);
and AND3 (N525, N522, N407, N215);
not NOT1 (N526, N503);
not NOT1 (N527, N525);
xor XOR2 (N528, N521, N92);
buf BUF1 (N529, N515);
xor XOR2 (N530, N518, N394);
buf BUF1 (N531, N493);
or OR3 (N532, N519, N317, N278);
xor XOR2 (N533, N531, N8);
buf BUF1 (N534, N495);
and AND4 (N535, N524, N382, N307, N89);
not NOT1 (N536, N530);
buf BUF1 (N537, N526);
xor XOR2 (N538, N523, N233);
not NOT1 (N539, N537);
not NOT1 (N540, N533);
or OR2 (N541, N540, N99);
xor XOR2 (N542, N539, N537);
and AND2 (N543, N528, N248);
xor XOR2 (N544, N534, N52);
nor NOR4 (N545, N532, N169, N106, N226);
nand NAND2 (N546, N542, N224);
buf BUF1 (N547, N541);
buf BUF1 (N548, N544);
buf BUF1 (N549, N527);
xor XOR2 (N550, N545, N352);
not NOT1 (N551, N529);
not NOT1 (N552, N543);
nor NOR3 (N553, N546, N87, N316);
xor XOR2 (N554, N548, N463);
buf BUF1 (N555, N553);
not NOT1 (N556, N538);
nand NAND4 (N557, N535, N475, N275, N18);
buf BUF1 (N558, N555);
xor XOR2 (N559, N558, N300);
nand NAND4 (N560, N559, N66, N268, N57);
or OR2 (N561, N551, N553);
and AND4 (N562, N547, N439, N175, N503);
buf BUF1 (N563, N552);
nand NAND2 (N564, N549, N294);
nor NOR3 (N565, N560, N204, N66);
or OR4 (N566, N565, N291, N242, N303);
xor XOR2 (N567, N561, N177);
xor XOR2 (N568, N567, N490);
or OR4 (N569, N563, N390, N358, N113);
and AND3 (N570, N569, N286, N330);
not NOT1 (N571, N568);
and AND3 (N572, N570, N254, N325);
buf BUF1 (N573, N556);
or OR2 (N574, N562, N39);
not NOT1 (N575, N566);
buf BUF1 (N576, N572);
buf BUF1 (N577, N550);
or OR3 (N578, N575, N87, N364);
and AND4 (N579, N564, N158, N452, N536);
and AND3 (N580, N517, N579, N180);
buf BUF1 (N581, N567);
xor XOR2 (N582, N578, N108);
not NOT1 (N583, N574);
nand NAND4 (N584, N571, N472, N261, N451);
nor NOR4 (N585, N554, N218, N552, N65);
or OR3 (N586, N581, N99, N287);
xor XOR2 (N587, N586, N569);
or OR4 (N588, N580, N400, N244, N362);
or OR3 (N589, N584, N15, N130);
buf BUF1 (N590, N589);
and AND3 (N591, N588, N14, N417);
and AND2 (N592, N590, N197);
nor NOR2 (N593, N577, N565);
nand NAND3 (N594, N593, N592, N65);
or OR3 (N595, N396, N161, N15);
xor XOR2 (N596, N557, N435);
not NOT1 (N597, N595);
xor XOR2 (N598, N583, N308);
or OR3 (N599, N598, N299, N158);
and AND2 (N600, N573, N259);
or OR2 (N601, N591, N204);
nor NOR3 (N602, N599, N534, N319);
xor XOR2 (N603, N585, N401);
nor NOR2 (N604, N602, N68);
buf BUF1 (N605, N603);
nand NAND2 (N606, N604, N161);
buf BUF1 (N607, N576);
xor XOR2 (N608, N601, N277);
xor XOR2 (N609, N600, N117);
and AND3 (N610, N582, N128, N233);
endmodule