// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;

output N8016,N8017,N8010,N8015,N7993,N8005,N8006,N8012,N7998,N8018;

nor NOR4 (N19, N14, N12, N10, N16);
nor NOR2 (N20, N8, N13);
not NOT1 (N21, N4);
buf BUF1 (N22, N12);
and AND3 (N23, N20, N13, N6);
xor XOR2 (N24, N12, N8);
or OR3 (N25, N21, N21, N18);
and AND3 (N26, N13, N23, N5);
nor NOR4 (N27, N14, N16, N13, N16);
xor XOR2 (N28, N12, N20);
not NOT1 (N29, N26);
nand NAND2 (N30, N17, N6);
and AND4 (N31, N3, N19, N10, N25);
nand NAND2 (N32, N31, N23);
not NOT1 (N33, N4);
nor NOR2 (N34, N11, N1);
buf BUF1 (N35, N16);
nor NOR3 (N36, N22, N5, N9);
xor XOR2 (N37, N32, N9);
nand NAND3 (N38, N36, N11, N35);
nand NAND3 (N39, N38, N34, N6);
not NOT1 (N40, N29);
buf BUF1 (N41, N14);
not NOT1 (N42, N25);
nand NAND3 (N43, N24, N15, N24);
not NOT1 (N44, N40);
not NOT1 (N45, N33);
and AND4 (N46, N37, N3, N16, N29);
nor NOR2 (N47, N41, N22);
not NOT1 (N48, N47);
and AND3 (N49, N27, N10, N15);
nor NOR2 (N50, N45, N32);
nand NAND4 (N51, N44, N48, N2, N22);
nand NAND2 (N52, N13, N40);
and AND2 (N53, N39, N47);
nor NOR2 (N54, N53, N7);
buf BUF1 (N55, N46);
nand NAND2 (N56, N42, N1);
and AND3 (N57, N50, N49, N53);
or OR2 (N58, N18, N35);
and AND3 (N59, N54, N41, N57);
not NOT1 (N60, N10);
and AND3 (N61, N55, N52, N37);
or OR3 (N62, N21, N39, N46);
and AND4 (N63, N59, N43, N53, N56);
nor NOR4 (N64, N29, N7, N59, N33);
xor XOR2 (N65, N13, N12);
xor XOR2 (N66, N51, N26);
not NOT1 (N67, N28);
nor NOR3 (N68, N60, N44, N58);
nand NAND4 (N69, N50, N23, N68, N45);
or OR4 (N70, N55, N52, N66, N64);
xor XOR2 (N71, N63, N54);
xor XOR2 (N72, N30, N31);
and AND2 (N73, N8, N23);
nor NOR4 (N74, N69, N48, N67, N11);
or OR4 (N75, N33, N45, N73, N50);
and AND3 (N76, N3, N57, N61);
not NOT1 (N77, N23);
not NOT1 (N78, N37);
nand NAND2 (N79, N74, N35);
nor NOR3 (N80, N75, N33, N31);
xor XOR2 (N81, N71, N48);
or OR3 (N82, N81, N77, N65);
nor NOR2 (N83, N27, N70);
xor XOR2 (N84, N26, N77);
buf BUF1 (N85, N76);
not NOT1 (N86, N13);
xor XOR2 (N87, N83, N49);
buf BUF1 (N88, N85);
nor NOR3 (N89, N72, N20, N19);
nor NOR3 (N90, N84, N63, N8);
not NOT1 (N91, N62);
buf BUF1 (N92, N87);
xor XOR2 (N93, N86, N16);
xor XOR2 (N94, N93, N2);
buf BUF1 (N95, N78);
nand NAND2 (N96, N92, N42);
nor NOR4 (N97, N91, N91, N75, N5);
and AND3 (N98, N90, N66, N29);
or OR2 (N99, N89, N64);
or OR4 (N100, N95, N87, N78, N52);
nor NOR3 (N101, N79, N7, N98);
nor NOR3 (N102, N38, N16, N66);
not NOT1 (N103, N97);
not NOT1 (N104, N99);
xor XOR2 (N105, N96, N79);
and AND3 (N106, N94, N15, N25);
nor NOR3 (N107, N103, N18, N82);
or OR2 (N108, N74, N63);
buf BUF1 (N109, N88);
not NOT1 (N110, N107);
and AND3 (N111, N101, N35, N70);
and AND2 (N112, N106, N102);
or OR4 (N113, N25, N47, N48, N86);
nand NAND4 (N114, N80, N6, N40, N26);
nand NAND3 (N115, N108, N114, N1);
and AND3 (N116, N41, N52, N78);
nor NOR2 (N117, N115, N38);
and AND4 (N118, N112, N74, N107, N75);
and AND4 (N119, N118, N96, N37, N37);
not NOT1 (N120, N116);
nand NAND3 (N121, N100, N25, N13);
xor XOR2 (N122, N111, N33);
nand NAND2 (N123, N110, N35);
not NOT1 (N124, N104);
not NOT1 (N125, N122);
not NOT1 (N126, N123);
or OR4 (N127, N119, N51, N86, N123);
nand NAND4 (N128, N125, N41, N24, N4);
and AND3 (N129, N128, N111, N123);
nand NAND3 (N130, N121, N110, N56);
xor XOR2 (N131, N113, N8);
and AND4 (N132, N124, N98, N95, N91);
nor NOR2 (N133, N126, N128);
nand NAND4 (N134, N130, N38, N122, N51);
or OR3 (N135, N105, N15, N82);
nor NOR2 (N136, N109, N26);
not NOT1 (N137, N129);
or OR4 (N138, N133, N41, N113, N108);
buf BUF1 (N139, N117);
and AND2 (N140, N138, N1);
not NOT1 (N141, N134);
xor XOR2 (N142, N141, N23);
xor XOR2 (N143, N139, N20);
buf BUF1 (N144, N135);
and AND2 (N145, N120, N131);
or OR3 (N146, N29, N61, N37);
and AND4 (N147, N127, N74, N17, N57);
xor XOR2 (N148, N132, N39);
buf BUF1 (N149, N147);
xor XOR2 (N150, N137, N71);
nor NOR3 (N151, N140, N125, N5);
xor XOR2 (N152, N149, N50);
or OR4 (N153, N145, N113, N2, N58);
nand NAND4 (N154, N136, N114, N107, N97);
not NOT1 (N155, N150);
and AND2 (N156, N152, N128);
buf BUF1 (N157, N146);
and AND2 (N158, N157, N6);
and AND4 (N159, N155, N57, N124, N61);
not NOT1 (N160, N142);
buf BUF1 (N161, N154);
not NOT1 (N162, N158);
buf BUF1 (N163, N144);
nand NAND3 (N164, N159, N73, N96);
xor XOR2 (N165, N148, N115);
not NOT1 (N166, N162);
and AND3 (N167, N153, N118, N128);
xor XOR2 (N168, N160, N78);
or OR2 (N169, N156, N42);
buf BUF1 (N170, N168);
nand NAND4 (N171, N151, N23, N30, N107);
xor XOR2 (N172, N171, N121);
not NOT1 (N173, N169);
xor XOR2 (N174, N172, N95);
and AND4 (N175, N143, N138, N15, N17);
nand NAND4 (N176, N163, N55, N32, N91);
or OR4 (N177, N174, N37, N110, N13);
buf BUF1 (N178, N166);
buf BUF1 (N179, N161);
nor NOR4 (N180, N178, N148, N168, N61);
xor XOR2 (N181, N173, N33);
nor NOR4 (N182, N164, N112, N70, N38);
nand NAND3 (N183, N180, N72, N26);
xor XOR2 (N184, N179, N82);
xor XOR2 (N185, N167, N45);
xor XOR2 (N186, N170, N60);
nor NOR3 (N187, N183, N167, N31);
and AND4 (N188, N176, N24, N93, N180);
xor XOR2 (N189, N182, N75);
xor XOR2 (N190, N184, N1);
nand NAND4 (N191, N165, N110, N62, N161);
and AND3 (N192, N188, N183, N105);
nand NAND2 (N193, N189, N155);
not NOT1 (N194, N187);
xor XOR2 (N195, N186, N133);
xor XOR2 (N196, N181, N16);
or OR4 (N197, N191, N193, N37, N68);
nand NAND2 (N198, N148, N197);
not NOT1 (N199, N97);
xor XOR2 (N200, N199, N13);
xor XOR2 (N201, N175, N100);
xor XOR2 (N202, N185, N145);
or OR3 (N203, N200, N202, N50);
nand NAND3 (N204, N175, N57, N13);
buf BUF1 (N205, N204);
xor XOR2 (N206, N205, N107);
nor NOR4 (N207, N203, N62, N197, N4);
xor XOR2 (N208, N190, N85);
nand NAND2 (N209, N206, N134);
buf BUF1 (N210, N208);
nand NAND2 (N211, N195, N68);
and AND2 (N212, N207, N121);
not NOT1 (N213, N198);
xor XOR2 (N214, N201, N100);
nand NAND3 (N215, N212, N114, N127);
buf BUF1 (N216, N215);
buf BUF1 (N217, N214);
nand NAND2 (N218, N216, N141);
buf BUF1 (N219, N192);
or OR4 (N220, N196, N202, N47, N7);
and AND2 (N221, N220, N147);
not NOT1 (N222, N209);
and AND2 (N223, N210, N215);
nor NOR3 (N224, N213, N188, N100);
or OR3 (N225, N223, N112, N155);
nand NAND2 (N226, N221, N21);
nor NOR3 (N227, N217, N169, N69);
and AND3 (N228, N225, N26, N85);
xor XOR2 (N229, N211, N196);
nand NAND4 (N230, N227, N40, N198, N66);
or OR3 (N231, N177, N142, N45);
nand NAND3 (N232, N224, N172, N206);
nor NOR3 (N233, N228, N96, N31);
nor NOR2 (N234, N218, N76);
nand NAND2 (N235, N232, N194);
not NOT1 (N236, N177);
nand NAND3 (N237, N233, N55, N17);
nor NOR4 (N238, N230, N5, N115, N44);
nand NAND2 (N239, N238, N88);
xor XOR2 (N240, N237, N137);
buf BUF1 (N241, N234);
not NOT1 (N242, N239);
nand NAND4 (N243, N240, N241, N148, N17);
or OR4 (N244, N192, N41, N30, N164);
or OR2 (N245, N236, N157);
buf BUF1 (N246, N235);
not NOT1 (N247, N226);
not NOT1 (N248, N219);
or OR2 (N249, N243, N151);
and AND3 (N250, N222, N130, N86);
or OR2 (N251, N229, N136);
nor NOR2 (N252, N250, N249);
buf BUF1 (N253, N25);
nor NOR2 (N254, N251, N206);
and AND3 (N255, N231, N121, N172);
nand NAND4 (N256, N252, N94, N209, N90);
not NOT1 (N257, N256);
buf BUF1 (N258, N245);
buf BUF1 (N259, N246);
nor NOR3 (N260, N247, N100, N14);
buf BUF1 (N261, N255);
nor NOR2 (N262, N253, N189);
nor NOR2 (N263, N244, N164);
nor NOR3 (N264, N257, N211, N140);
not NOT1 (N265, N263);
not NOT1 (N266, N264);
or OR4 (N267, N259, N251, N87, N163);
not NOT1 (N268, N258);
and AND4 (N269, N267, N51, N175, N131);
not NOT1 (N270, N269);
xor XOR2 (N271, N254, N71);
or OR2 (N272, N248, N215);
nor NOR4 (N273, N260, N107, N73, N16);
nand NAND4 (N274, N270, N160, N124, N72);
buf BUF1 (N275, N272);
or OR2 (N276, N274, N179);
or OR2 (N277, N273, N34);
or OR2 (N278, N261, N54);
and AND4 (N279, N268, N244, N160, N102);
not NOT1 (N280, N265);
xor XOR2 (N281, N278, N218);
nor NOR3 (N282, N279, N54, N82);
nor NOR3 (N283, N276, N177, N1);
nand NAND4 (N284, N262, N139, N8, N91);
xor XOR2 (N285, N266, N38);
nand NAND3 (N286, N275, N193, N242);
nand NAND4 (N287, N215, N101, N190, N126);
xor XOR2 (N288, N281, N103);
and AND3 (N289, N286, N250, N128);
nor NOR2 (N290, N288, N163);
nand NAND2 (N291, N271, N273);
buf BUF1 (N292, N289);
not NOT1 (N293, N284);
nand NAND3 (N294, N285, N177, N68);
nand NAND2 (N295, N294, N67);
not NOT1 (N296, N290);
or OR4 (N297, N283, N188, N280, N17);
not NOT1 (N298, N94);
nor NOR4 (N299, N298, N38, N279, N95);
nor NOR2 (N300, N297, N45);
xor XOR2 (N301, N287, N68);
or OR2 (N302, N296, N132);
not NOT1 (N303, N299);
nand NAND2 (N304, N301, N165);
nand NAND2 (N305, N293, N29);
buf BUF1 (N306, N291);
or OR2 (N307, N305, N121);
or OR2 (N308, N295, N110);
nand NAND2 (N309, N303, N24);
or OR4 (N310, N300, N73, N230, N64);
nand NAND3 (N311, N307, N242, N5);
or OR2 (N312, N302, N291);
and AND3 (N313, N304, N173, N219);
nor NOR3 (N314, N308, N124, N82);
or OR4 (N315, N310, N188, N83, N142);
nand NAND4 (N316, N277, N267, N122, N83);
xor XOR2 (N317, N315, N232);
buf BUF1 (N318, N292);
nand NAND2 (N319, N318, N205);
not NOT1 (N320, N319);
xor XOR2 (N321, N309, N46);
or OR4 (N322, N316, N300, N318, N180);
nor NOR4 (N323, N306, N312, N31, N265);
nor NOR2 (N324, N225, N201);
nand NAND4 (N325, N324, N302, N285, N194);
xor XOR2 (N326, N282, N95);
xor XOR2 (N327, N323, N119);
not NOT1 (N328, N325);
xor XOR2 (N329, N314, N7);
xor XOR2 (N330, N311, N115);
and AND2 (N331, N320, N40);
not NOT1 (N332, N327);
xor XOR2 (N333, N317, N216);
nor NOR2 (N334, N331, N328);
or OR2 (N335, N266, N203);
buf BUF1 (N336, N329);
nor NOR4 (N337, N335, N117, N186, N79);
buf BUF1 (N338, N322);
and AND3 (N339, N334, N122, N305);
not NOT1 (N340, N339);
xor XOR2 (N341, N313, N13);
xor XOR2 (N342, N336, N45);
or OR4 (N343, N333, N209, N222, N21);
nor NOR3 (N344, N321, N213, N92);
xor XOR2 (N345, N344, N114);
buf BUF1 (N346, N342);
not NOT1 (N347, N332);
or OR4 (N348, N341, N105, N299, N309);
buf BUF1 (N349, N330);
nor NOR3 (N350, N347, N339, N187);
nand NAND2 (N351, N338, N69);
and AND2 (N352, N348, N24);
xor XOR2 (N353, N345, N212);
not NOT1 (N354, N351);
buf BUF1 (N355, N349);
xor XOR2 (N356, N326, N259);
nor NOR3 (N357, N340, N29, N65);
nor NOR3 (N358, N352, N134, N336);
and AND2 (N359, N353, N311);
not NOT1 (N360, N359);
nor NOR2 (N361, N350, N199);
nand NAND2 (N362, N346, N226);
and AND2 (N363, N360, N26);
buf BUF1 (N364, N363);
or OR2 (N365, N354, N57);
not NOT1 (N366, N355);
not NOT1 (N367, N365);
buf BUF1 (N368, N362);
nand NAND3 (N369, N358, N294, N321);
nor NOR3 (N370, N356, N104, N130);
nand NAND2 (N371, N369, N137);
or OR2 (N372, N371, N283);
nor NOR2 (N373, N366, N116);
nor NOR3 (N374, N337, N281, N271);
and AND3 (N375, N367, N157, N67);
buf BUF1 (N376, N368);
and AND3 (N377, N343, N320, N325);
or OR4 (N378, N375, N33, N177, N129);
and AND4 (N379, N364, N212, N93, N148);
and AND4 (N380, N378, N142, N301, N158);
xor XOR2 (N381, N377, N318);
buf BUF1 (N382, N381);
nor NOR2 (N383, N361, N22);
not NOT1 (N384, N376);
nor NOR2 (N385, N373, N278);
nor NOR2 (N386, N380, N21);
not NOT1 (N387, N374);
or OR2 (N388, N383, N315);
nor NOR2 (N389, N384, N237);
nand NAND4 (N390, N379, N76, N382, N120);
buf BUF1 (N391, N253);
or OR4 (N392, N370, N153, N154, N287);
not NOT1 (N393, N386);
nand NAND2 (N394, N389, N2);
nand NAND3 (N395, N372, N164, N183);
not NOT1 (N396, N388);
xor XOR2 (N397, N390, N329);
and AND3 (N398, N357, N310, N218);
or OR2 (N399, N392, N331);
not NOT1 (N400, N399);
nand NAND4 (N401, N396, N337, N363, N145);
nor NOR2 (N402, N401, N327);
and AND4 (N403, N393, N24, N302, N16);
or OR2 (N404, N391, N40);
nor NOR4 (N405, N402, N316, N171, N181);
buf BUF1 (N406, N404);
not NOT1 (N407, N398);
and AND2 (N408, N406, N42);
buf BUF1 (N409, N405);
xor XOR2 (N410, N407, N150);
or OR2 (N411, N408, N234);
nor NOR4 (N412, N411, N41, N276, N132);
nand NAND4 (N413, N385, N82, N208, N216);
buf BUF1 (N414, N413);
or OR4 (N415, N403, N166, N56, N288);
xor XOR2 (N416, N400, N135);
or OR4 (N417, N394, N70, N213, N172);
nand NAND4 (N418, N410, N127, N328, N268);
nand NAND4 (N419, N414, N56, N91, N159);
nor NOR4 (N420, N397, N136, N102, N85);
nand NAND4 (N421, N418, N241, N365, N286);
buf BUF1 (N422, N420);
buf BUF1 (N423, N395);
xor XOR2 (N424, N412, N336);
nor NOR4 (N425, N424, N411, N198, N378);
not NOT1 (N426, N387);
not NOT1 (N427, N422);
nor NOR4 (N428, N423, N23, N185, N170);
nand NAND4 (N429, N421, N114, N11, N219);
xor XOR2 (N430, N415, N339);
or OR2 (N431, N430, N72);
nand NAND2 (N432, N425, N389);
xor XOR2 (N433, N427, N48);
nor NOR3 (N434, N433, N316, N47);
buf BUF1 (N435, N429);
nor NOR3 (N436, N426, N128, N141);
buf BUF1 (N437, N416);
buf BUF1 (N438, N428);
buf BUF1 (N439, N432);
not NOT1 (N440, N409);
or OR4 (N441, N417, N360, N235, N350);
buf BUF1 (N442, N437);
not NOT1 (N443, N435);
or OR2 (N444, N441, N202);
nor NOR3 (N445, N436, N201, N84);
and AND2 (N446, N442, N219);
buf BUF1 (N447, N440);
and AND2 (N448, N431, N222);
nor NOR3 (N449, N434, N99, N402);
and AND3 (N450, N444, N317, N105);
nand NAND4 (N451, N438, N130, N390, N243);
not NOT1 (N452, N448);
nor NOR3 (N453, N451, N197, N374);
nor NOR2 (N454, N419, N219);
buf BUF1 (N455, N453);
or OR3 (N456, N439, N109, N17);
and AND2 (N457, N454, N202);
or OR4 (N458, N452, N193, N444, N36);
nor NOR2 (N459, N458, N380);
or OR3 (N460, N459, N100, N53);
buf BUF1 (N461, N447);
or OR4 (N462, N450, N66, N417, N409);
or OR3 (N463, N446, N317, N428);
nor NOR3 (N464, N445, N327, N305);
and AND4 (N465, N464, N422, N424, N265);
nor NOR2 (N466, N443, N394);
not NOT1 (N467, N462);
buf BUF1 (N468, N467);
not NOT1 (N469, N456);
xor XOR2 (N470, N457, N226);
buf BUF1 (N471, N455);
or OR4 (N472, N469, N443, N30, N26);
or OR4 (N473, N463, N222, N369, N334);
nand NAND3 (N474, N449, N26, N28);
and AND4 (N475, N465, N171, N324, N2);
nor NOR2 (N476, N461, N430);
nand NAND3 (N477, N466, N347, N46);
nor NOR3 (N478, N473, N468, N360);
buf BUF1 (N479, N246);
buf BUF1 (N480, N472);
not NOT1 (N481, N471);
nor NOR2 (N482, N470, N234);
nor NOR3 (N483, N460, N383, N51);
xor XOR2 (N484, N480, N324);
or OR2 (N485, N477, N344);
or OR2 (N486, N476, N108);
buf BUF1 (N487, N484);
buf BUF1 (N488, N481);
or OR3 (N489, N483, N21, N285);
xor XOR2 (N490, N488, N83);
and AND4 (N491, N486, N112, N24, N367);
nor NOR2 (N492, N479, N141);
and AND2 (N493, N475, N372);
and AND3 (N494, N490, N222, N258);
buf BUF1 (N495, N492);
nor NOR2 (N496, N474, N189);
not NOT1 (N497, N495);
not NOT1 (N498, N493);
nor NOR2 (N499, N478, N425);
xor XOR2 (N500, N485, N460);
or OR3 (N501, N496, N51, N381);
buf BUF1 (N502, N489);
xor XOR2 (N503, N497, N203);
or OR4 (N504, N498, N454, N104, N202);
or OR2 (N505, N502, N91);
or OR4 (N506, N499, N400, N383, N500);
buf BUF1 (N507, N50);
or OR4 (N508, N501, N32, N200, N169);
or OR2 (N509, N503, N181);
nor NOR2 (N510, N506, N223);
or OR3 (N511, N508, N94, N473);
nor NOR4 (N512, N482, N151, N255, N226);
or OR3 (N513, N487, N206, N416);
and AND2 (N514, N494, N364);
buf BUF1 (N515, N514);
xor XOR2 (N516, N512, N192);
nand NAND2 (N517, N515, N51);
nand NAND4 (N518, N507, N319, N98, N381);
and AND3 (N519, N491, N312, N444);
buf BUF1 (N520, N504);
not NOT1 (N521, N517);
xor XOR2 (N522, N505, N34);
xor XOR2 (N523, N522, N288);
not NOT1 (N524, N519);
not NOT1 (N525, N523);
xor XOR2 (N526, N525, N400);
nand NAND3 (N527, N526, N406, N101);
and AND2 (N528, N521, N173);
xor XOR2 (N529, N524, N401);
xor XOR2 (N530, N511, N43);
xor XOR2 (N531, N510, N278);
xor XOR2 (N532, N527, N311);
not NOT1 (N533, N513);
nor NOR3 (N534, N532, N412, N252);
and AND2 (N535, N529, N109);
nand NAND4 (N536, N520, N138, N490, N249);
buf BUF1 (N537, N535);
xor XOR2 (N538, N531, N32);
xor XOR2 (N539, N536, N160);
nor NOR2 (N540, N534, N388);
buf BUF1 (N541, N539);
xor XOR2 (N542, N530, N466);
and AND4 (N543, N509, N275, N165, N2);
or OR4 (N544, N528, N373, N363, N373);
xor XOR2 (N545, N516, N226);
buf BUF1 (N546, N544);
nand NAND4 (N547, N518, N494, N287, N264);
nand NAND4 (N548, N533, N416, N359, N91);
or OR2 (N549, N538, N229);
or OR2 (N550, N548, N426);
not NOT1 (N551, N549);
buf BUF1 (N552, N541);
buf BUF1 (N553, N537);
nor NOR4 (N554, N553, N300, N241, N65);
or OR4 (N555, N552, N330, N554, N208);
or OR3 (N556, N106, N401, N71);
and AND3 (N557, N550, N322, N363);
nor NOR2 (N558, N556, N242);
nand NAND3 (N559, N546, N120, N281);
or OR3 (N560, N543, N14, N204);
nand NAND2 (N561, N557, N296);
not NOT1 (N562, N540);
nor NOR3 (N563, N558, N520, N327);
nor NOR3 (N564, N542, N370, N153);
xor XOR2 (N565, N562, N120);
not NOT1 (N566, N547);
not NOT1 (N567, N561);
or OR3 (N568, N564, N5, N97);
buf BUF1 (N569, N567);
xor XOR2 (N570, N551, N559);
nand NAND4 (N571, N416, N377, N387, N94);
and AND3 (N572, N565, N207, N120);
xor XOR2 (N573, N563, N282);
or OR2 (N574, N568, N256);
nand NAND2 (N575, N572, N427);
nor NOR3 (N576, N570, N449, N261);
buf BUF1 (N577, N545);
buf BUF1 (N578, N576);
xor XOR2 (N579, N571, N100);
nand NAND4 (N580, N575, N516, N152, N561);
not NOT1 (N581, N573);
nor NOR3 (N582, N578, N36, N515);
buf BUF1 (N583, N560);
xor XOR2 (N584, N580, N73);
and AND4 (N585, N577, N557, N114, N576);
buf BUF1 (N586, N585);
nand NAND4 (N587, N579, N357, N569, N171);
or OR4 (N588, N24, N52, N17, N460);
nor NOR3 (N589, N555, N506, N57);
buf BUF1 (N590, N587);
buf BUF1 (N591, N590);
not NOT1 (N592, N581);
xor XOR2 (N593, N582, N501);
nor NOR2 (N594, N586, N327);
not NOT1 (N595, N566);
buf BUF1 (N596, N591);
buf BUF1 (N597, N592);
not NOT1 (N598, N584);
and AND4 (N599, N596, N362, N243, N394);
nor NOR3 (N600, N593, N225, N587);
or OR2 (N601, N588, N580);
nor NOR2 (N602, N589, N346);
buf BUF1 (N603, N602);
or OR2 (N604, N599, N453);
or OR3 (N605, N598, N494, N475);
xor XOR2 (N606, N594, N570);
xor XOR2 (N607, N600, N138);
or OR3 (N608, N604, N328, N398);
not NOT1 (N609, N608);
nor NOR2 (N610, N574, N199);
nor NOR2 (N611, N605, N495);
xor XOR2 (N612, N610, N352);
xor XOR2 (N613, N595, N483);
nand NAND2 (N614, N609, N289);
and AND4 (N615, N603, N71, N315, N461);
nor NOR4 (N616, N597, N311, N53, N291);
xor XOR2 (N617, N616, N144);
nor NOR3 (N618, N607, N116, N381);
nand NAND4 (N619, N583, N240, N296, N198);
or OR4 (N620, N619, N304, N459, N583);
or OR2 (N621, N611, N431);
xor XOR2 (N622, N606, N441);
and AND2 (N623, N613, N187);
buf BUF1 (N624, N617);
xor XOR2 (N625, N615, N589);
and AND4 (N626, N622, N420, N30, N324);
or OR4 (N627, N601, N344, N204, N453);
xor XOR2 (N628, N612, N597);
or OR4 (N629, N625, N168, N442, N5);
and AND3 (N630, N621, N151, N548);
buf BUF1 (N631, N624);
nor NOR3 (N632, N630, N185, N177);
and AND4 (N633, N620, N557, N293, N231);
and AND3 (N634, N632, N404, N307);
not NOT1 (N635, N618);
buf BUF1 (N636, N633);
buf BUF1 (N637, N631);
nor NOR2 (N638, N628, N19);
or OR2 (N639, N627, N380);
not NOT1 (N640, N629);
nand NAND2 (N641, N634, N539);
buf BUF1 (N642, N635);
buf BUF1 (N643, N639);
or OR3 (N644, N641, N107, N444);
nor NOR2 (N645, N623, N576);
nand NAND4 (N646, N642, N515, N43, N258);
or OR4 (N647, N638, N15, N368, N482);
nor NOR3 (N648, N645, N605, N497);
xor XOR2 (N649, N626, N334);
xor XOR2 (N650, N636, N229);
nand NAND2 (N651, N643, N310);
xor XOR2 (N652, N648, N291);
not NOT1 (N653, N637);
and AND3 (N654, N647, N220, N377);
xor XOR2 (N655, N646, N387);
not NOT1 (N656, N652);
xor XOR2 (N657, N653, N39);
nand NAND2 (N658, N656, N154);
and AND3 (N659, N640, N536, N114);
and AND4 (N660, N657, N63, N278, N260);
buf BUF1 (N661, N650);
xor XOR2 (N662, N649, N487);
not NOT1 (N663, N660);
not NOT1 (N664, N662);
xor XOR2 (N665, N664, N22);
buf BUF1 (N666, N651);
not NOT1 (N667, N665);
or OR4 (N668, N614, N551, N127, N340);
xor XOR2 (N669, N668, N245);
and AND2 (N670, N666, N121);
nand NAND2 (N671, N659, N627);
not NOT1 (N672, N667);
buf BUF1 (N673, N661);
nand NAND2 (N674, N672, N489);
nor NOR2 (N675, N658, N56);
and AND4 (N676, N670, N263, N19, N503);
nand NAND3 (N677, N644, N672, N661);
xor XOR2 (N678, N675, N106);
xor XOR2 (N679, N673, N42);
not NOT1 (N680, N663);
nand NAND4 (N681, N674, N537, N287, N394);
nand NAND2 (N682, N679, N550);
buf BUF1 (N683, N655);
or OR4 (N684, N681, N491, N541, N503);
and AND3 (N685, N680, N668, N161);
nor NOR2 (N686, N682, N401);
buf BUF1 (N687, N678);
or OR2 (N688, N687, N237);
nand NAND2 (N689, N677, N140);
not NOT1 (N690, N683);
and AND2 (N691, N689, N344);
nand NAND4 (N692, N690, N602, N21, N308);
buf BUF1 (N693, N691);
nor NOR3 (N694, N669, N225, N139);
xor XOR2 (N695, N671, N54);
nor NOR2 (N696, N695, N243);
nand NAND3 (N697, N676, N115, N25);
and AND4 (N698, N684, N659, N235, N57);
or OR4 (N699, N696, N398, N105, N31);
not NOT1 (N700, N686);
xor XOR2 (N701, N698, N696);
buf BUF1 (N702, N688);
xor XOR2 (N703, N693, N571);
nand NAND3 (N704, N701, N23, N425);
and AND4 (N705, N694, N407, N485, N609);
buf BUF1 (N706, N685);
and AND2 (N707, N700, N355);
buf BUF1 (N708, N702);
buf BUF1 (N709, N707);
nor NOR4 (N710, N706, N199, N79, N620);
xor XOR2 (N711, N709, N505);
or OR3 (N712, N692, N599, N69);
nor NOR2 (N713, N697, N14);
xor XOR2 (N714, N704, N98);
buf BUF1 (N715, N699);
nand NAND3 (N716, N705, N163, N488);
xor XOR2 (N717, N710, N424);
and AND2 (N718, N654, N190);
nand NAND3 (N719, N713, N664, N625);
not NOT1 (N720, N719);
nand NAND3 (N721, N715, N490, N716);
not NOT1 (N722, N431);
nand NAND3 (N723, N703, N201, N282);
nor NOR2 (N724, N718, N599);
nand NAND2 (N725, N714, N713);
not NOT1 (N726, N720);
and AND4 (N727, N725, N209, N103, N614);
buf BUF1 (N728, N726);
or OR4 (N729, N724, N392, N678, N236);
and AND2 (N730, N728, N146);
buf BUF1 (N731, N729);
buf BUF1 (N732, N723);
xor XOR2 (N733, N708, N575);
nor NOR3 (N734, N711, N189, N46);
and AND3 (N735, N722, N352, N286);
xor XOR2 (N736, N730, N203);
xor XOR2 (N737, N735, N695);
xor XOR2 (N738, N712, N208);
nand NAND4 (N739, N738, N553, N185, N172);
nand NAND3 (N740, N727, N141, N587);
nand NAND2 (N741, N717, N555);
and AND3 (N742, N736, N159, N241);
and AND3 (N743, N742, N435, N476);
xor XOR2 (N744, N721, N35);
nand NAND3 (N745, N733, N683, N431);
buf BUF1 (N746, N743);
or OR3 (N747, N744, N742, N254);
nand NAND3 (N748, N745, N531, N171);
buf BUF1 (N749, N747);
xor XOR2 (N750, N746, N109);
nand NAND3 (N751, N732, N421, N366);
and AND3 (N752, N750, N301, N601);
xor XOR2 (N753, N731, N266);
not NOT1 (N754, N751);
nand NAND4 (N755, N734, N640, N578, N138);
buf BUF1 (N756, N739);
not NOT1 (N757, N740);
nor NOR3 (N758, N737, N268, N248);
not NOT1 (N759, N752);
not NOT1 (N760, N756);
nand NAND2 (N761, N749, N396);
xor XOR2 (N762, N753, N9);
nor NOR2 (N763, N755, N91);
and AND2 (N764, N757, N315);
xor XOR2 (N765, N760, N558);
nand NAND2 (N766, N754, N330);
or OR4 (N767, N761, N354, N219, N508);
nor NOR4 (N768, N748, N164, N148, N736);
not NOT1 (N769, N765);
and AND2 (N770, N769, N366);
not NOT1 (N771, N767);
nand NAND2 (N772, N768, N24);
nor NOR4 (N773, N771, N424, N238, N416);
nor NOR2 (N774, N762, N124);
not NOT1 (N775, N758);
nor NOR2 (N776, N741, N479);
and AND4 (N777, N773, N229, N743, N599);
nand NAND4 (N778, N774, N597, N298, N308);
not NOT1 (N779, N777);
xor XOR2 (N780, N759, N640);
nor NOR3 (N781, N766, N270, N86);
or OR2 (N782, N770, N321);
nor NOR2 (N783, N764, N357);
not NOT1 (N784, N778);
and AND3 (N785, N763, N781, N560);
and AND3 (N786, N175, N239, N686);
xor XOR2 (N787, N772, N167);
xor XOR2 (N788, N780, N564);
nor NOR3 (N789, N786, N175, N366);
or OR3 (N790, N787, N648, N305);
or OR4 (N791, N775, N332, N773, N572);
and AND3 (N792, N784, N554, N432);
nand NAND3 (N793, N783, N94, N615);
nor NOR4 (N794, N793, N271, N81, N185);
buf BUF1 (N795, N782);
nor NOR2 (N796, N789, N329);
xor XOR2 (N797, N776, N337);
xor XOR2 (N798, N797, N210);
nand NAND3 (N799, N779, N334, N515);
or OR3 (N800, N799, N761, N221);
or OR3 (N801, N795, N716, N575);
or OR2 (N802, N791, N29);
nand NAND2 (N803, N798, N548);
buf BUF1 (N804, N796);
or OR3 (N805, N794, N498, N485);
or OR3 (N806, N792, N508, N538);
nor NOR4 (N807, N802, N91, N179, N443);
nor NOR2 (N808, N801, N307);
not NOT1 (N809, N804);
and AND4 (N810, N807, N211, N355, N593);
buf BUF1 (N811, N785);
nand NAND2 (N812, N808, N685);
nand NAND4 (N813, N812, N201, N530, N204);
xor XOR2 (N814, N810, N62);
and AND3 (N815, N800, N602, N428);
nand NAND3 (N816, N813, N267, N187);
xor XOR2 (N817, N816, N164);
buf BUF1 (N818, N806);
nand NAND2 (N819, N818, N464);
buf BUF1 (N820, N805);
and AND4 (N821, N814, N812, N285, N57);
nor NOR4 (N822, N809, N535, N37, N248);
nand NAND2 (N823, N821, N730);
nand NAND2 (N824, N819, N536);
and AND3 (N825, N823, N132, N806);
buf BUF1 (N826, N788);
buf BUF1 (N827, N811);
and AND3 (N828, N824, N394, N477);
buf BUF1 (N829, N790);
or OR4 (N830, N820, N205, N111, N181);
xor XOR2 (N831, N827, N115);
or OR4 (N832, N822, N224, N782, N649);
or OR4 (N833, N829, N378, N120, N201);
and AND2 (N834, N817, N278);
not NOT1 (N835, N828);
and AND4 (N836, N833, N496, N628, N50);
nand NAND2 (N837, N826, N461);
nand NAND3 (N838, N815, N174, N688);
nand NAND2 (N839, N836, N808);
nand NAND2 (N840, N839, N42);
not NOT1 (N841, N831);
or OR4 (N842, N841, N617, N419, N219);
and AND4 (N843, N835, N205, N52, N395);
or OR2 (N844, N837, N554);
nor NOR3 (N845, N825, N536, N370);
nor NOR3 (N846, N838, N780, N324);
or OR2 (N847, N843, N511);
nand NAND2 (N848, N847, N229);
buf BUF1 (N849, N832);
xor XOR2 (N850, N845, N740);
and AND4 (N851, N803, N387, N745, N826);
not NOT1 (N852, N840);
or OR4 (N853, N846, N78, N403, N620);
xor XOR2 (N854, N850, N241);
buf BUF1 (N855, N849);
not NOT1 (N856, N834);
nand NAND2 (N857, N844, N147);
xor XOR2 (N858, N848, N809);
xor XOR2 (N859, N858, N117);
or OR4 (N860, N842, N264, N511, N378);
nor NOR4 (N861, N830, N517, N1, N649);
buf BUF1 (N862, N852);
nand NAND4 (N863, N851, N215, N98, N22);
nand NAND2 (N864, N856, N359);
xor XOR2 (N865, N854, N161);
nand NAND3 (N866, N859, N212, N700);
xor XOR2 (N867, N853, N537);
nand NAND4 (N868, N867, N323, N791, N558);
xor XOR2 (N869, N855, N99);
xor XOR2 (N870, N868, N4);
buf BUF1 (N871, N865);
not NOT1 (N872, N862);
not NOT1 (N873, N871);
nor NOR3 (N874, N873, N871, N790);
buf BUF1 (N875, N863);
or OR2 (N876, N864, N386);
not NOT1 (N877, N869);
not NOT1 (N878, N866);
or OR4 (N879, N877, N155, N608, N7);
xor XOR2 (N880, N872, N522);
not NOT1 (N881, N861);
buf BUF1 (N882, N876);
not NOT1 (N883, N857);
or OR2 (N884, N870, N74);
nand NAND2 (N885, N860, N336);
or OR2 (N886, N878, N32);
buf BUF1 (N887, N881);
xor XOR2 (N888, N875, N596);
nor NOR4 (N889, N886, N459, N494, N630);
or OR2 (N890, N888, N412);
nand NAND2 (N891, N885, N334);
and AND2 (N892, N879, N802);
xor XOR2 (N893, N887, N618);
nor NOR2 (N894, N882, N790);
nand NAND2 (N895, N894, N297);
or OR2 (N896, N895, N432);
nor NOR4 (N897, N896, N774, N222, N321);
nor NOR3 (N898, N891, N384, N518);
not NOT1 (N899, N880);
not NOT1 (N900, N899);
buf BUF1 (N901, N889);
not NOT1 (N902, N890);
and AND4 (N903, N897, N170, N857, N124);
nor NOR3 (N904, N901, N3, N681);
nor NOR2 (N905, N892, N388);
not NOT1 (N906, N900);
nor NOR2 (N907, N884, N20);
not NOT1 (N908, N902);
not NOT1 (N909, N906);
and AND2 (N910, N907, N868);
or OR2 (N911, N905, N888);
or OR2 (N912, N908, N861);
nor NOR4 (N913, N911, N581, N558, N513);
xor XOR2 (N914, N883, N175);
not NOT1 (N915, N904);
nor NOR4 (N916, N874, N84, N187, N715);
buf BUF1 (N917, N913);
nor NOR2 (N918, N912, N434);
or OR4 (N919, N898, N563, N583, N624);
not NOT1 (N920, N918);
xor XOR2 (N921, N903, N866);
or OR4 (N922, N919, N563, N535, N410);
and AND2 (N923, N910, N263);
nor NOR4 (N924, N917, N452, N302, N431);
nand NAND2 (N925, N923, N519);
or OR4 (N926, N920, N643, N719, N360);
and AND2 (N927, N926, N259);
and AND4 (N928, N924, N241, N775, N534);
nor NOR4 (N929, N914, N841, N543, N530);
not NOT1 (N930, N909);
and AND3 (N931, N915, N69, N762);
xor XOR2 (N932, N930, N608);
and AND3 (N933, N931, N500, N637);
or OR3 (N934, N925, N902, N125);
and AND2 (N935, N928, N290);
not NOT1 (N936, N932);
buf BUF1 (N937, N933);
not NOT1 (N938, N893);
buf BUF1 (N939, N938);
nor NOR2 (N940, N927, N579);
buf BUF1 (N941, N940);
nand NAND2 (N942, N936, N553);
or OR4 (N943, N934, N704, N370, N121);
xor XOR2 (N944, N937, N508);
or OR3 (N945, N942, N428, N96);
or OR3 (N946, N939, N741, N94);
and AND3 (N947, N945, N871, N555);
not NOT1 (N948, N947);
buf BUF1 (N949, N941);
xor XOR2 (N950, N948, N932);
nor NOR3 (N951, N950, N848, N290);
or OR2 (N952, N921, N669);
and AND2 (N953, N951, N699);
not NOT1 (N954, N922);
buf BUF1 (N955, N943);
xor XOR2 (N956, N952, N197);
nor NOR3 (N957, N953, N914, N428);
or OR4 (N958, N944, N498, N716, N209);
or OR3 (N959, N946, N416, N79);
xor XOR2 (N960, N957, N667);
or OR2 (N961, N955, N348);
nand NAND3 (N962, N929, N305, N715);
nor NOR2 (N963, N956, N151);
nor NOR2 (N964, N961, N613);
nand NAND4 (N965, N962, N474, N829, N538);
or OR4 (N966, N965, N623, N175, N274);
nor NOR3 (N967, N964, N455, N59);
not NOT1 (N968, N960);
xor XOR2 (N969, N963, N450);
xor XOR2 (N970, N949, N482);
nor NOR3 (N971, N935, N790, N630);
buf BUF1 (N972, N916);
buf BUF1 (N973, N967);
not NOT1 (N974, N968);
nand NAND3 (N975, N973, N486, N367);
not NOT1 (N976, N958);
buf BUF1 (N977, N954);
buf BUF1 (N978, N977);
buf BUF1 (N979, N976);
not NOT1 (N980, N979);
xor XOR2 (N981, N969, N186);
xor XOR2 (N982, N980, N247);
or OR3 (N983, N974, N701, N800);
nor NOR2 (N984, N981, N803);
nor NOR2 (N985, N982, N258);
not NOT1 (N986, N971);
xor XOR2 (N987, N986, N507);
not NOT1 (N988, N972);
xor XOR2 (N989, N985, N388);
xor XOR2 (N990, N978, N327);
nor NOR4 (N991, N990, N672, N40, N2);
xor XOR2 (N992, N989, N555);
nor NOR4 (N993, N984, N598, N12, N464);
nor NOR3 (N994, N975, N320, N916);
xor XOR2 (N995, N966, N917);
xor XOR2 (N996, N991, N956);
xor XOR2 (N997, N970, N787);
and AND4 (N998, N959, N942, N556, N867);
xor XOR2 (N999, N988, N837);
xor XOR2 (N1000, N996, N997);
and AND2 (N1001, N701, N144);
xor XOR2 (N1002, N987, N396);
nand NAND3 (N1003, N999, N819, N631);
or OR2 (N1004, N1000, N594);
not NOT1 (N1005, N998);
and AND3 (N1006, N994, N336, N912);
nor NOR2 (N1007, N993, N747);
or OR4 (N1008, N983, N489, N896, N75);
buf BUF1 (N1009, N1008);
and AND2 (N1010, N1001, N475);
xor XOR2 (N1011, N1005, N662);
and AND3 (N1012, N1004, N729, N839);
nand NAND3 (N1013, N1002, N642, N739);
or OR2 (N1014, N1009, N683);
nand NAND3 (N1015, N1007, N872, N16);
or OR2 (N1016, N1010, N612);
nand NAND3 (N1017, N995, N788, N31);
nor NOR4 (N1018, N1015, N498, N307, N69);
buf BUF1 (N1019, N1011);
not NOT1 (N1020, N1019);
xor XOR2 (N1021, N1014, N186);
not NOT1 (N1022, N1012);
buf BUF1 (N1023, N1006);
and AND3 (N1024, N1013, N483, N857);
xor XOR2 (N1025, N1016, N105);
or OR2 (N1026, N1022, N630);
xor XOR2 (N1027, N1003, N167);
or OR3 (N1028, N1020, N759, N621);
and AND2 (N1029, N1018, N163);
and AND4 (N1030, N1028, N747, N198, N306);
nand NAND2 (N1031, N1024, N799);
or OR2 (N1032, N992, N578);
nor NOR4 (N1033, N1025, N67, N251, N325);
or OR4 (N1034, N1033, N425, N847, N622);
buf BUF1 (N1035, N1023);
buf BUF1 (N1036, N1032);
and AND4 (N1037, N1030, N371, N77, N16);
nor NOR2 (N1038, N1031, N575);
buf BUF1 (N1039, N1021);
or OR4 (N1040, N1017, N446, N288, N989);
or OR2 (N1041, N1036, N607);
and AND4 (N1042, N1035, N201, N850, N760);
not NOT1 (N1043, N1040);
nor NOR4 (N1044, N1039, N254, N983, N985);
not NOT1 (N1045, N1044);
xor XOR2 (N1046, N1043, N692);
nor NOR3 (N1047, N1041, N90, N429);
nor NOR3 (N1048, N1029, N127, N10);
and AND4 (N1049, N1026, N965, N704, N925);
nand NAND3 (N1050, N1045, N1041, N59);
not NOT1 (N1051, N1038);
and AND3 (N1052, N1046, N20, N514);
buf BUF1 (N1053, N1027);
not NOT1 (N1054, N1050);
or OR2 (N1055, N1052, N521);
and AND4 (N1056, N1042, N272, N334, N739);
nand NAND4 (N1057, N1056, N842, N574, N266);
not NOT1 (N1058, N1051);
and AND3 (N1059, N1037, N734, N395);
not NOT1 (N1060, N1057);
xor XOR2 (N1061, N1055, N165);
not NOT1 (N1062, N1053);
and AND4 (N1063, N1062, N437, N922, N26);
buf BUF1 (N1064, N1063);
not NOT1 (N1065, N1047);
buf BUF1 (N1066, N1054);
xor XOR2 (N1067, N1058, N973);
or OR2 (N1068, N1064, N480);
xor XOR2 (N1069, N1065, N547);
nand NAND2 (N1070, N1067, N713);
buf BUF1 (N1071, N1060);
nand NAND4 (N1072, N1068, N457, N598, N307);
nand NAND4 (N1073, N1061, N914, N391, N520);
xor XOR2 (N1074, N1049, N21);
and AND4 (N1075, N1048, N235, N451, N960);
buf BUF1 (N1076, N1066);
xor XOR2 (N1077, N1069, N849);
buf BUF1 (N1078, N1059);
nor NOR2 (N1079, N1073, N871);
nor NOR3 (N1080, N1079, N241, N147);
nand NAND3 (N1081, N1072, N764, N605);
and AND4 (N1082, N1080, N123, N859, N76);
buf BUF1 (N1083, N1034);
or OR4 (N1084, N1081, N102, N1038, N299);
nand NAND2 (N1085, N1082, N131);
or OR4 (N1086, N1071, N976, N204, N56);
and AND3 (N1087, N1070, N859, N916);
buf BUF1 (N1088, N1077);
and AND3 (N1089, N1075, N175, N1073);
buf BUF1 (N1090, N1089);
nor NOR2 (N1091, N1090, N1063);
not NOT1 (N1092, N1086);
nand NAND4 (N1093, N1087, N760, N367, N541);
nor NOR3 (N1094, N1092, N572, N606);
xor XOR2 (N1095, N1083, N890);
nor NOR3 (N1096, N1074, N551, N72);
and AND3 (N1097, N1096, N7, N272);
xor XOR2 (N1098, N1078, N127);
nor NOR4 (N1099, N1084, N460, N216, N899);
buf BUF1 (N1100, N1094);
xor XOR2 (N1101, N1099, N278);
nand NAND3 (N1102, N1101, N862, N542);
buf BUF1 (N1103, N1102);
or OR4 (N1104, N1076, N584, N827, N708);
nand NAND4 (N1105, N1091, N822, N429, N130);
and AND4 (N1106, N1100, N614, N949, N790);
not NOT1 (N1107, N1093);
xor XOR2 (N1108, N1103, N391);
buf BUF1 (N1109, N1098);
not NOT1 (N1110, N1088);
and AND3 (N1111, N1097, N904, N663);
xor XOR2 (N1112, N1106, N995);
or OR2 (N1113, N1104, N861);
nand NAND2 (N1114, N1112, N151);
nor NOR4 (N1115, N1108, N967, N1082, N78);
nand NAND3 (N1116, N1105, N253, N1066);
or OR2 (N1117, N1113, N996);
xor XOR2 (N1118, N1114, N761);
or OR3 (N1119, N1117, N457, N1058);
or OR3 (N1120, N1116, N106, N608);
xor XOR2 (N1121, N1095, N436);
nand NAND3 (N1122, N1119, N6, N1104);
buf BUF1 (N1123, N1121);
buf BUF1 (N1124, N1110);
buf BUF1 (N1125, N1109);
nand NAND3 (N1126, N1107, N121, N734);
buf BUF1 (N1127, N1085);
nand NAND2 (N1128, N1122, N834);
not NOT1 (N1129, N1125);
not NOT1 (N1130, N1127);
and AND4 (N1131, N1120, N620, N46, N1053);
or OR2 (N1132, N1124, N485);
nand NAND4 (N1133, N1123, N837, N290, N507);
and AND3 (N1134, N1131, N17, N420);
nand NAND4 (N1135, N1133, N593, N245, N605);
nand NAND2 (N1136, N1111, N583);
xor XOR2 (N1137, N1134, N266);
nor NOR4 (N1138, N1129, N793, N203, N586);
not NOT1 (N1139, N1135);
or OR3 (N1140, N1118, N652, N690);
or OR4 (N1141, N1137, N28, N607, N403);
or OR4 (N1142, N1136, N834, N913, N462);
not NOT1 (N1143, N1141);
nor NOR3 (N1144, N1139, N101, N314);
xor XOR2 (N1145, N1128, N221);
xor XOR2 (N1146, N1144, N617);
nand NAND4 (N1147, N1142, N806, N476, N884);
and AND4 (N1148, N1132, N527, N745, N241);
buf BUF1 (N1149, N1140);
not NOT1 (N1150, N1138);
nor NOR4 (N1151, N1148, N132, N259, N49);
buf BUF1 (N1152, N1151);
nand NAND2 (N1153, N1152, N1073);
nand NAND3 (N1154, N1153, N686, N75);
nor NOR4 (N1155, N1150, N492, N153, N227);
buf BUF1 (N1156, N1130);
nand NAND4 (N1157, N1149, N957, N329, N636);
xor XOR2 (N1158, N1157, N128);
buf BUF1 (N1159, N1147);
and AND4 (N1160, N1156, N151, N430, N505);
nand NAND3 (N1161, N1143, N528, N169);
nor NOR3 (N1162, N1155, N187, N1095);
nor NOR4 (N1163, N1162, N632, N180, N508);
nand NAND2 (N1164, N1158, N772);
and AND4 (N1165, N1126, N889, N1135, N452);
xor XOR2 (N1166, N1163, N894);
buf BUF1 (N1167, N1166);
and AND2 (N1168, N1160, N893);
nor NOR4 (N1169, N1145, N331, N698, N119);
not NOT1 (N1170, N1164);
xor XOR2 (N1171, N1146, N10);
nand NAND2 (N1172, N1170, N769);
and AND3 (N1173, N1169, N1125, N486);
or OR3 (N1174, N1172, N546, N1172);
buf BUF1 (N1175, N1159);
not NOT1 (N1176, N1168);
nand NAND4 (N1177, N1176, N764, N761, N243);
not NOT1 (N1178, N1165);
not NOT1 (N1179, N1115);
nor NOR2 (N1180, N1179, N730);
or OR4 (N1181, N1171, N976, N565, N1100);
or OR3 (N1182, N1154, N493, N845);
nand NAND2 (N1183, N1161, N694);
and AND3 (N1184, N1167, N1058, N988);
and AND2 (N1185, N1175, N141);
and AND3 (N1186, N1180, N284, N838);
buf BUF1 (N1187, N1173);
and AND2 (N1188, N1184, N41);
xor XOR2 (N1189, N1188, N787);
xor XOR2 (N1190, N1189, N458);
buf BUF1 (N1191, N1185);
nand NAND3 (N1192, N1181, N955, N921);
not NOT1 (N1193, N1178);
buf BUF1 (N1194, N1186);
buf BUF1 (N1195, N1193);
not NOT1 (N1196, N1174);
and AND2 (N1197, N1183, N759);
not NOT1 (N1198, N1191);
buf BUF1 (N1199, N1195);
xor XOR2 (N1200, N1187, N272);
buf BUF1 (N1201, N1198);
buf BUF1 (N1202, N1177);
not NOT1 (N1203, N1201);
nand NAND4 (N1204, N1197, N319, N393, N658);
xor XOR2 (N1205, N1182, N1045);
and AND2 (N1206, N1192, N708);
nand NAND2 (N1207, N1190, N1086);
xor XOR2 (N1208, N1202, N614);
nand NAND4 (N1209, N1206, N29, N156, N678);
not NOT1 (N1210, N1203);
not NOT1 (N1211, N1196);
nor NOR4 (N1212, N1208, N387, N22, N124);
buf BUF1 (N1213, N1210);
xor XOR2 (N1214, N1194, N1034);
nand NAND3 (N1215, N1200, N970, N359);
or OR2 (N1216, N1213, N483);
or OR2 (N1217, N1205, N1021);
and AND3 (N1218, N1214, N185, N227);
buf BUF1 (N1219, N1207);
buf BUF1 (N1220, N1215);
nor NOR2 (N1221, N1211, N1078);
or OR4 (N1222, N1199, N285, N117, N626);
or OR4 (N1223, N1212, N115, N293, N766);
xor XOR2 (N1224, N1223, N1015);
xor XOR2 (N1225, N1204, N667);
nand NAND2 (N1226, N1225, N360);
not NOT1 (N1227, N1220);
or OR2 (N1228, N1226, N871);
nand NAND3 (N1229, N1209, N822, N1194);
nand NAND2 (N1230, N1222, N1199);
buf BUF1 (N1231, N1224);
nand NAND3 (N1232, N1229, N1117, N551);
or OR3 (N1233, N1231, N773, N1039);
or OR3 (N1234, N1219, N85, N918);
and AND2 (N1235, N1227, N566);
and AND3 (N1236, N1217, N708, N518);
nor NOR2 (N1237, N1234, N1175);
not NOT1 (N1238, N1235);
buf BUF1 (N1239, N1236);
xor XOR2 (N1240, N1238, N364);
buf BUF1 (N1241, N1218);
or OR2 (N1242, N1228, N242);
not NOT1 (N1243, N1237);
xor XOR2 (N1244, N1216, N1);
buf BUF1 (N1245, N1221);
nand NAND3 (N1246, N1244, N562, N272);
nor NOR2 (N1247, N1233, N1105);
nand NAND2 (N1248, N1246, N651);
not NOT1 (N1249, N1230);
not NOT1 (N1250, N1241);
nand NAND2 (N1251, N1248, N1035);
and AND4 (N1252, N1243, N34, N551, N798);
or OR2 (N1253, N1247, N626);
or OR2 (N1254, N1251, N438);
not NOT1 (N1255, N1254);
buf BUF1 (N1256, N1252);
nand NAND4 (N1257, N1240, N931, N1169, N633);
xor XOR2 (N1258, N1245, N972);
buf BUF1 (N1259, N1232);
nor NOR4 (N1260, N1249, N405, N158, N388);
or OR4 (N1261, N1255, N127, N1182, N634);
not NOT1 (N1262, N1242);
buf BUF1 (N1263, N1253);
nor NOR2 (N1264, N1262, N279);
buf BUF1 (N1265, N1260);
or OR2 (N1266, N1239, N261);
xor XOR2 (N1267, N1257, N385);
buf BUF1 (N1268, N1259);
xor XOR2 (N1269, N1261, N327);
nand NAND3 (N1270, N1256, N874, N622);
not NOT1 (N1271, N1263);
or OR2 (N1272, N1250, N992);
and AND4 (N1273, N1269, N1231, N345, N380);
nand NAND4 (N1274, N1265, N403, N443, N796);
nor NOR4 (N1275, N1267, N138, N453, N190);
xor XOR2 (N1276, N1270, N1091);
nand NAND2 (N1277, N1275, N461);
nor NOR3 (N1278, N1274, N88, N577);
buf BUF1 (N1279, N1278);
xor XOR2 (N1280, N1258, N507);
and AND2 (N1281, N1277, N1206);
and AND4 (N1282, N1271, N1201, N1137, N43);
and AND3 (N1283, N1281, N599, N828);
not NOT1 (N1284, N1280);
xor XOR2 (N1285, N1268, N145);
not NOT1 (N1286, N1282);
and AND4 (N1287, N1286, N1091, N489, N201);
buf BUF1 (N1288, N1272);
buf BUF1 (N1289, N1266);
and AND3 (N1290, N1288, N509, N84);
and AND4 (N1291, N1273, N15, N981, N526);
not NOT1 (N1292, N1285);
nand NAND4 (N1293, N1264, N1286, N267, N339);
xor XOR2 (N1294, N1291, N490);
and AND2 (N1295, N1289, N374);
or OR2 (N1296, N1290, N808);
or OR2 (N1297, N1294, N536);
nand NAND3 (N1298, N1292, N138, N576);
nand NAND2 (N1299, N1283, N930);
nand NAND2 (N1300, N1297, N611);
and AND4 (N1301, N1293, N1006, N1055, N613);
and AND2 (N1302, N1300, N1161);
or OR4 (N1303, N1301, N202, N1118, N345);
and AND4 (N1304, N1296, N834, N132, N742);
nand NAND2 (N1305, N1304, N631);
nand NAND4 (N1306, N1295, N652, N838, N398);
nor NOR4 (N1307, N1284, N788, N891, N617);
or OR4 (N1308, N1287, N462, N59, N697);
nand NAND2 (N1309, N1306, N162);
nand NAND2 (N1310, N1307, N669);
buf BUF1 (N1311, N1310);
xor XOR2 (N1312, N1276, N1188);
or OR3 (N1313, N1312, N1009, N874);
buf BUF1 (N1314, N1302);
xor XOR2 (N1315, N1279, N1240);
or OR4 (N1316, N1313, N282, N1054, N676);
nor NOR4 (N1317, N1308, N527, N995, N116);
nor NOR2 (N1318, N1317, N981);
buf BUF1 (N1319, N1316);
buf BUF1 (N1320, N1314);
nor NOR3 (N1321, N1299, N773, N863);
xor XOR2 (N1322, N1318, N1243);
or OR4 (N1323, N1309, N273, N545, N191);
nor NOR4 (N1324, N1315, N238, N989, N1189);
nand NAND2 (N1325, N1303, N211);
and AND4 (N1326, N1319, N1112, N867, N373);
nor NOR2 (N1327, N1311, N5);
buf BUF1 (N1328, N1323);
nor NOR2 (N1329, N1321, N124);
xor XOR2 (N1330, N1322, N953);
or OR4 (N1331, N1324, N1296, N46, N1186);
not NOT1 (N1332, N1298);
not NOT1 (N1333, N1329);
not NOT1 (N1334, N1305);
xor XOR2 (N1335, N1325, N1279);
nand NAND4 (N1336, N1328, N165, N778, N35);
and AND2 (N1337, N1335, N962);
nor NOR3 (N1338, N1320, N1018, N871);
nor NOR3 (N1339, N1326, N235, N523);
and AND3 (N1340, N1333, N324, N981);
xor XOR2 (N1341, N1330, N741);
and AND3 (N1342, N1337, N1192, N995);
not NOT1 (N1343, N1336);
nor NOR4 (N1344, N1341, N1257, N1164, N612);
xor XOR2 (N1345, N1342, N348);
and AND2 (N1346, N1345, N33);
xor XOR2 (N1347, N1339, N67);
xor XOR2 (N1348, N1327, N1212);
and AND4 (N1349, N1346, N1133, N737, N88);
nor NOR4 (N1350, N1334, N294, N841, N213);
not NOT1 (N1351, N1343);
nand NAND3 (N1352, N1331, N1252, N963);
not NOT1 (N1353, N1338);
or OR3 (N1354, N1344, N710, N358);
not NOT1 (N1355, N1351);
not NOT1 (N1356, N1340);
buf BUF1 (N1357, N1355);
and AND4 (N1358, N1350, N624, N1256, N966);
buf BUF1 (N1359, N1348);
and AND4 (N1360, N1356, N104, N125, N340);
and AND4 (N1361, N1360, N161, N165, N264);
buf BUF1 (N1362, N1353);
not NOT1 (N1363, N1362);
nand NAND2 (N1364, N1352, N296);
xor XOR2 (N1365, N1358, N370);
buf BUF1 (N1366, N1364);
and AND4 (N1367, N1361, N49, N1096, N667);
xor XOR2 (N1368, N1349, N1354);
nand NAND2 (N1369, N719, N157);
buf BUF1 (N1370, N1368);
or OR2 (N1371, N1367, N603);
or OR4 (N1372, N1359, N573, N522, N1143);
and AND3 (N1373, N1372, N335, N990);
xor XOR2 (N1374, N1373, N101);
not NOT1 (N1375, N1347);
nor NOR2 (N1376, N1363, N1186);
xor XOR2 (N1377, N1332, N646);
not NOT1 (N1378, N1365);
xor XOR2 (N1379, N1374, N894);
nor NOR2 (N1380, N1378, N411);
nor NOR2 (N1381, N1379, N1093);
not NOT1 (N1382, N1371);
xor XOR2 (N1383, N1370, N1075);
and AND2 (N1384, N1369, N1332);
xor XOR2 (N1385, N1377, N882);
buf BUF1 (N1386, N1385);
not NOT1 (N1387, N1376);
buf BUF1 (N1388, N1387);
and AND3 (N1389, N1386, N925, N1182);
nor NOR4 (N1390, N1380, N806, N657, N908);
nor NOR2 (N1391, N1382, N63);
nand NAND2 (N1392, N1390, N988);
nand NAND4 (N1393, N1391, N439, N232, N972);
and AND3 (N1394, N1381, N744, N238);
xor XOR2 (N1395, N1384, N904);
nand NAND2 (N1396, N1393, N495);
nor NOR3 (N1397, N1383, N538, N625);
nor NOR3 (N1398, N1357, N329, N200);
or OR2 (N1399, N1388, N702);
nand NAND3 (N1400, N1392, N717, N707);
buf BUF1 (N1401, N1397);
and AND2 (N1402, N1400, N1032);
and AND2 (N1403, N1401, N672);
xor XOR2 (N1404, N1394, N114);
nand NAND2 (N1405, N1375, N833);
not NOT1 (N1406, N1404);
xor XOR2 (N1407, N1399, N499);
xor XOR2 (N1408, N1366, N804);
and AND3 (N1409, N1389, N1349, N334);
not NOT1 (N1410, N1395);
xor XOR2 (N1411, N1407, N62);
xor XOR2 (N1412, N1405, N1387);
xor XOR2 (N1413, N1409, N457);
not NOT1 (N1414, N1413);
nand NAND4 (N1415, N1411, N1354, N647, N1293);
buf BUF1 (N1416, N1406);
xor XOR2 (N1417, N1416, N224);
nor NOR3 (N1418, N1408, N281, N903);
and AND4 (N1419, N1412, N60, N653, N624);
not NOT1 (N1420, N1398);
nor NOR3 (N1421, N1415, N1288, N460);
nand NAND2 (N1422, N1418, N162);
nand NAND4 (N1423, N1421, N1057, N684, N192);
xor XOR2 (N1424, N1410, N509);
and AND2 (N1425, N1396, N1357);
nand NAND4 (N1426, N1423, N1168, N688, N520);
buf BUF1 (N1427, N1403);
buf BUF1 (N1428, N1425);
xor XOR2 (N1429, N1402, N760);
xor XOR2 (N1430, N1422, N347);
buf BUF1 (N1431, N1417);
buf BUF1 (N1432, N1420);
or OR4 (N1433, N1414, N551, N866, N575);
nand NAND3 (N1434, N1424, N26, N939);
nand NAND2 (N1435, N1419, N1256);
and AND4 (N1436, N1435, N152, N1423, N1092);
not NOT1 (N1437, N1431);
and AND3 (N1438, N1434, N994, N1231);
or OR4 (N1439, N1438, N543, N491, N1155);
xor XOR2 (N1440, N1437, N1068);
not NOT1 (N1441, N1432);
or OR2 (N1442, N1429, N1124);
xor XOR2 (N1443, N1428, N242);
xor XOR2 (N1444, N1433, N409);
or OR4 (N1445, N1444, N643, N1000, N809);
and AND2 (N1446, N1440, N1264);
buf BUF1 (N1447, N1446);
nor NOR3 (N1448, N1447, N843, N163);
xor XOR2 (N1449, N1443, N504);
xor XOR2 (N1450, N1449, N308);
and AND2 (N1451, N1442, N940);
or OR4 (N1452, N1451, N748, N4, N39);
buf BUF1 (N1453, N1450);
not NOT1 (N1454, N1426);
nand NAND3 (N1455, N1441, N1168, N252);
and AND4 (N1456, N1427, N241, N861, N8);
or OR3 (N1457, N1436, N102, N284);
and AND2 (N1458, N1452, N591);
and AND4 (N1459, N1430, N682, N1283, N384);
and AND2 (N1460, N1459, N1341);
or OR3 (N1461, N1455, N455, N1411);
xor XOR2 (N1462, N1448, N975);
xor XOR2 (N1463, N1458, N150);
nand NAND4 (N1464, N1462, N578, N1142, N289);
and AND3 (N1465, N1453, N614, N238);
not NOT1 (N1466, N1460);
buf BUF1 (N1467, N1465);
or OR2 (N1468, N1454, N127);
buf BUF1 (N1469, N1466);
and AND4 (N1470, N1467, N1148, N897, N626);
nor NOR4 (N1471, N1457, N1116, N667, N1234);
xor XOR2 (N1472, N1469, N82);
buf BUF1 (N1473, N1470);
buf BUF1 (N1474, N1472);
or OR2 (N1475, N1463, N392);
xor XOR2 (N1476, N1464, N604);
or OR4 (N1477, N1468, N857, N1423, N1259);
not NOT1 (N1478, N1476);
not NOT1 (N1479, N1478);
not NOT1 (N1480, N1477);
xor XOR2 (N1481, N1480, N1446);
nor NOR4 (N1482, N1461, N302, N911, N780);
not NOT1 (N1483, N1473);
not NOT1 (N1484, N1456);
not NOT1 (N1485, N1475);
nor NOR4 (N1486, N1483, N763, N172, N1475);
or OR2 (N1487, N1471, N1339);
xor XOR2 (N1488, N1439, N127);
and AND2 (N1489, N1474, N977);
nand NAND2 (N1490, N1489, N76);
and AND3 (N1491, N1445, N433, N172);
or OR2 (N1492, N1482, N898);
or OR2 (N1493, N1486, N102);
nand NAND4 (N1494, N1493, N386, N422, N1065);
or OR4 (N1495, N1479, N838, N242, N1033);
or OR2 (N1496, N1490, N537);
nand NAND3 (N1497, N1481, N596, N842);
or OR3 (N1498, N1497, N1446, N1315);
nand NAND2 (N1499, N1491, N803);
nor NOR3 (N1500, N1487, N1123, N309);
nor NOR4 (N1501, N1498, N980, N15, N375);
buf BUF1 (N1502, N1496);
or OR3 (N1503, N1499, N1452, N1009);
buf BUF1 (N1504, N1500);
nor NOR4 (N1505, N1504, N883, N1287, N1220);
or OR4 (N1506, N1488, N312, N1337, N235);
xor XOR2 (N1507, N1494, N742);
and AND3 (N1508, N1505, N62, N1480);
nand NAND3 (N1509, N1485, N653, N1248);
nand NAND3 (N1510, N1503, N630, N746);
nand NAND2 (N1511, N1509, N707);
xor XOR2 (N1512, N1492, N1021);
or OR4 (N1513, N1484, N227, N815, N77);
xor XOR2 (N1514, N1512, N914);
xor XOR2 (N1515, N1506, N665);
nand NAND2 (N1516, N1515, N316);
and AND4 (N1517, N1516, N314, N1035, N1065);
xor XOR2 (N1518, N1495, N127);
buf BUF1 (N1519, N1511);
or OR4 (N1520, N1514, N202, N549, N273);
not NOT1 (N1521, N1513);
or OR4 (N1522, N1518, N1068, N753, N1477);
nand NAND4 (N1523, N1501, N77, N28, N699);
buf BUF1 (N1524, N1522);
and AND4 (N1525, N1519, N1403, N638, N416);
not NOT1 (N1526, N1507);
nor NOR4 (N1527, N1525, N130, N746, N811);
or OR4 (N1528, N1526, N956, N1174, N1227);
xor XOR2 (N1529, N1508, N1442);
nor NOR4 (N1530, N1521, N753, N1373, N1178);
or OR4 (N1531, N1528, N96, N1078, N475);
buf BUF1 (N1532, N1510);
not NOT1 (N1533, N1520);
xor XOR2 (N1534, N1532, N909);
or OR4 (N1535, N1527, N606, N1041, N1373);
and AND4 (N1536, N1530, N1227, N415, N850);
nand NAND2 (N1537, N1534, N322);
buf BUF1 (N1538, N1537);
buf BUF1 (N1539, N1524);
and AND3 (N1540, N1539, N586, N1493);
nor NOR4 (N1541, N1533, N1190, N849, N197);
nor NOR2 (N1542, N1536, N766);
nand NAND3 (N1543, N1523, N573, N805);
nand NAND4 (N1544, N1540, N1030, N1079, N60);
buf BUF1 (N1545, N1542);
nor NOR3 (N1546, N1535, N1027, N920);
nor NOR2 (N1547, N1546, N1481);
or OR2 (N1548, N1541, N1171);
nand NAND2 (N1549, N1538, N1032);
buf BUF1 (N1550, N1545);
or OR2 (N1551, N1547, N1380);
or OR4 (N1552, N1529, N1484, N1259, N543);
nand NAND4 (N1553, N1548, N927, N234, N1280);
xor XOR2 (N1554, N1543, N281);
and AND4 (N1555, N1550, N623, N230, N1076);
and AND2 (N1556, N1554, N1090);
and AND2 (N1557, N1556, N605);
nand NAND2 (N1558, N1557, N990);
nand NAND3 (N1559, N1549, N68, N190);
nor NOR4 (N1560, N1517, N887, N255, N11);
xor XOR2 (N1561, N1560, N831);
or OR4 (N1562, N1555, N889, N20, N63);
nor NOR4 (N1563, N1552, N918, N1282, N708);
xor XOR2 (N1564, N1553, N746);
nor NOR4 (N1565, N1531, N158, N75, N1267);
xor XOR2 (N1566, N1565, N605);
buf BUF1 (N1567, N1551);
buf BUF1 (N1568, N1559);
buf BUF1 (N1569, N1558);
buf BUF1 (N1570, N1563);
nor NOR3 (N1571, N1544, N146, N4);
nor NOR2 (N1572, N1571, N1296);
buf BUF1 (N1573, N1562);
not NOT1 (N1574, N1566);
nor NOR2 (N1575, N1569, N457);
nor NOR2 (N1576, N1572, N1121);
xor XOR2 (N1577, N1561, N913);
or OR3 (N1578, N1570, N840, N454);
and AND2 (N1579, N1502, N1362);
nand NAND4 (N1580, N1574, N1282, N1133, N167);
not NOT1 (N1581, N1575);
and AND3 (N1582, N1577, N251, N712);
or OR3 (N1583, N1582, N1441, N1148);
or OR2 (N1584, N1578, N1407);
not NOT1 (N1585, N1568);
not NOT1 (N1586, N1583);
not NOT1 (N1587, N1567);
or OR2 (N1588, N1573, N812);
or OR4 (N1589, N1579, N1094, N1085, N1276);
not NOT1 (N1590, N1581);
buf BUF1 (N1591, N1576);
or OR2 (N1592, N1587, N29);
and AND2 (N1593, N1585, N781);
nor NOR2 (N1594, N1592, N1294);
xor XOR2 (N1595, N1589, N598);
nor NOR3 (N1596, N1586, N39, N285);
buf BUF1 (N1597, N1595);
buf BUF1 (N1598, N1588);
nand NAND3 (N1599, N1584, N1116, N132);
nor NOR3 (N1600, N1590, N1260, N1088);
nor NOR3 (N1601, N1593, N100, N1542);
buf BUF1 (N1602, N1598);
xor XOR2 (N1603, N1591, N394);
nand NAND4 (N1604, N1594, N368, N1206, N1400);
buf BUF1 (N1605, N1604);
and AND2 (N1606, N1597, N471);
xor XOR2 (N1607, N1600, N447);
and AND3 (N1608, N1599, N1581, N1480);
xor XOR2 (N1609, N1607, N798);
nand NAND3 (N1610, N1564, N1171, N211);
or OR3 (N1611, N1580, N762, N1596);
or OR2 (N1612, N638, N1177);
nor NOR2 (N1613, N1609, N1257);
nor NOR2 (N1614, N1606, N75);
nor NOR3 (N1615, N1601, N855, N1274);
and AND3 (N1616, N1615, N1322, N422);
nand NAND4 (N1617, N1602, N882, N679, N537);
nand NAND4 (N1618, N1613, N138, N862, N1404);
or OR2 (N1619, N1618, N909);
xor XOR2 (N1620, N1610, N998);
or OR2 (N1621, N1617, N1564);
nor NOR4 (N1622, N1620, N386, N161, N243);
nand NAND2 (N1623, N1611, N1296);
nand NAND3 (N1624, N1614, N3, N1575);
nor NOR2 (N1625, N1622, N153);
not NOT1 (N1626, N1608);
not NOT1 (N1627, N1625);
not NOT1 (N1628, N1616);
xor XOR2 (N1629, N1603, N115);
buf BUF1 (N1630, N1605);
or OR2 (N1631, N1630, N213);
buf BUF1 (N1632, N1612);
xor XOR2 (N1633, N1632, N1260);
nor NOR4 (N1634, N1629, N255, N610, N590);
and AND3 (N1635, N1633, N44, N194);
or OR3 (N1636, N1634, N1175, N1306);
xor XOR2 (N1637, N1627, N922);
nor NOR3 (N1638, N1631, N918, N60);
or OR2 (N1639, N1626, N1615);
nand NAND4 (N1640, N1621, N521, N370, N316);
nor NOR4 (N1641, N1639, N1207, N495, N724);
nand NAND3 (N1642, N1623, N174, N570);
nor NOR3 (N1643, N1638, N778, N1343);
nand NAND4 (N1644, N1635, N803, N1199, N1593);
not NOT1 (N1645, N1641);
xor XOR2 (N1646, N1628, N1224);
not NOT1 (N1647, N1645);
buf BUF1 (N1648, N1647);
nand NAND3 (N1649, N1636, N81, N1551);
xor XOR2 (N1650, N1619, N138);
nor NOR4 (N1651, N1650, N1404, N882, N138);
nand NAND2 (N1652, N1646, N470);
buf BUF1 (N1653, N1644);
nor NOR2 (N1654, N1637, N1532);
not NOT1 (N1655, N1653);
or OR2 (N1656, N1655, N419);
xor XOR2 (N1657, N1648, N1585);
xor XOR2 (N1658, N1640, N1272);
xor XOR2 (N1659, N1624, N297);
buf BUF1 (N1660, N1642);
nand NAND2 (N1661, N1652, N1439);
not NOT1 (N1662, N1659);
or OR3 (N1663, N1657, N345, N1451);
or OR4 (N1664, N1643, N630, N295, N1347);
not NOT1 (N1665, N1656);
or OR3 (N1666, N1660, N817, N440);
buf BUF1 (N1667, N1665);
xor XOR2 (N1668, N1661, N1535);
nand NAND2 (N1669, N1664, N982);
xor XOR2 (N1670, N1669, N1294);
or OR2 (N1671, N1666, N175);
nor NOR2 (N1672, N1662, N772);
buf BUF1 (N1673, N1663);
nor NOR4 (N1674, N1658, N875, N1021, N113);
nor NOR4 (N1675, N1671, N995, N523, N418);
or OR3 (N1676, N1672, N1119, N241);
not NOT1 (N1677, N1667);
and AND4 (N1678, N1675, N137, N1148, N831);
or OR2 (N1679, N1676, N1294);
and AND4 (N1680, N1668, N27, N237, N668);
and AND2 (N1681, N1680, N1344);
xor XOR2 (N1682, N1677, N1619);
xor XOR2 (N1683, N1678, N336);
nor NOR2 (N1684, N1674, N1662);
not NOT1 (N1685, N1679);
nor NOR2 (N1686, N1670, N1646);
nand NAND2 (N1687, N1673, N1015);
and AND2 (N1688, N1685, N774);
not NOT1 (N1689, N1681);
nor NOR2 (N1690, N1651, N209);
and AND2 (N1691, N1682, N382);
nor NOR2 (N1692, N1654, N739);
or OR3 (N1693, N1692, N258, N1011);
nor NOR3 (N1694, N1684, N1219, N1687);
not NOT1 (N1695, N1461);
nor NOR3 (N1696, N1688, N1395, N875);
nor NOR4 (N1697, N1695, N492, N987, N1560);
or OR3 (N1698, N1649, N1665, N476);
buf BUF1 (N1699, N1683);
buf BUF1 (N1700, N1696);
buf BUF1 (N1701, N1686);
nor NOR3 (N1702, N1697, N935, N147);
nor NOR3 (N1703, N1699, N911, N286);
nor NOR3 (N1704, N1694, N66, N647);
nor NOR3 (N1705, N1702, N1135, N1440);
and AND2 (N1706, N1693, N71);
xor XOR2 (N1707, N1701, N1206);
nand NAND2 (N1708, N1691, N684);
xor XOR2 (N1709, N1700, N1240);
and AND4 (N1710, N1709, N934, N568, N677);
or OR4 (N1711, N1698, N1090, N1175, N1671);
or OR3 (N1712, N1690, N1476, N608);
xor XOR2 (N1713, N1689, N1114);
buf BUF1 (N1714, N1713);
buf BUF1 (N1715, N1704);
nand NAND2 (N1716, N1708, N802);
and AND3 (N1717, N1705, N285, N317);
xor XOR2 (N1718, N1711, N607);
xor XOR2 (N1719, N1703, N1463);
buf BUF1 (N1720, N1718);
nand NAND3 (N1721, N1719, N1447, N711);
buf BUF1 (N1722, N1716);
nor NOR2 (N1723, N1720, N647);
and AND4 (N1724, N1722, N1166, N1628, N1170);
and AND2 (N1725, N1712, N1250);
buf BUF1 (N1726, N1706);
nand NAND2 (N1727, N1725, N1534);
nor NOR2 (N1728, N1717, N1663);
buf BUF1 (N1729, N1707);
or OR2 (N1730, N1714, N172);
nor NOR3 (N1731, N1728, N926, N852);
nand NAND2 (N1732, N1729, N1366);
or OR4 (N1733, N1731, N1050, N1292, N1428);
or OR3 (N1734, N1724, N1356, N1129);
not NOT1 (N1735, N1730);
nor NOR3 (N1736, N1715, N875, N1457);
not NOT1 (N1737, N1710);
nor NOR2 (N1738, N1735, N1001);
nand NAND4 (N1739, N1727, N70, N435, N483);
xor XOR2 (N1740, N1721, N524);
and AND2 (N1741, N1734, N142);
nand NAND4 (N1742, N1739, N382, N177, N936);
nor NOR4 (N1743, N1726, N777, N1471, N292);
buf BUF1 (N1744, N1732);
and AND3 (N1745, N1723, N1447, N1242);
xor XOR2 (N1746, N1740, N1660);
or OR3 (N1747, N1733, N1742, N891);
and AND3 (N1748, N1454, N782, N1213);
nor NOR3 (N1749, N1743, N542, N315);
xor XOR2 (N1750, N1748, N191);
or OR3 (N1751, N1747, N1725, N465);
buf BUF1 (N1752, N1741);
buf BUF1 (N1753, N1752);
xor XOR2 (N1754, N1744, N355);
nand NAND4 (N1755, N1745, N1334, N953, N1688);
buf BUF1 (N1756, N1746);
buf BUF1 (N1757, N1751);
nor NOR4 (N1758, N1750, N1297, N203, N375);
xor XOR2 (N1759, N1758, N1246);
and AND3 (N1760, N1738, N1738, N1263);
and AND2 (N1761, N1753, N504);
and AND2 (N1762, N1757, N595);
buf BUF1 (N1763, N1759);
nand NAND4 (N1764, N1756, N1088, N1591, N341);
xor XOR2 (N1765, N1737, N188);
nor NOR2 (N1766, N1765, N405);
nor NOR3 (N1767, N1755, N751, N1433);
and AND4 (N1768, N1767, N134, N219, N1438);
or OR4 (N1769, N1749, N910, N182, N1153);
or OR2 (N1770, N1763, N1158);
or OR4 (N1771, N1736, N1451, N62, N742);
nand NAND4 (N1772, N1764, N1130, N664, N663);
and AND3 (N1773, N1760, N968, N1616);
not NOT1 (N1774, N1762);
nand NAND3 (N1775, N1761, N656, N1565);
xor XOR2 (N1776, N1772, N823);
xor XOR2 (N1777, N1773, N1147);
nand NAND2 (N1778, N1766, N614);
nor NOR2 (N1779, N1771, N838);
xor XOR2 (N1780, N1777, N115);
xor XOR2 (N1781, N1776, N84);
buf BUF1 (N1782, N1781);
and AND2 (N1783, N1775, N1542);
not NOT1 (N1784, N1754);
and AND4 (N1785, N1782, N935, N1060, N1066);
nor NOR2 (N1786, N1780, N294);
nor NOR2 (N1787, N1784, N1446);
not NOT1 (N1788, N1774);
nor NOR4 (N1789, N1779, N217, N704, N1379);
not NOT1 (N1790, N1778);
and AND4 (N1791, N1789, N878, N784, N750);
and AND2 (N1792, N1770, N732);
buf BUF1 (N1793, N1785);
not NOT1 (N1794, N1792);
xor XOR2 (N1795, N1768, N1168);
nand NAND3 (N1796, N1791, N1592, N714);
not NOT1 (N1797, N1795);
or OR2 (N1798, N1793, N21);
or OR3 (N1799, N1769, N1103, N1302);
buf BUF1 (N1800, N1790);
nand NAND4 (N1801, N1794, N1654, N1641, N196);
or OR4 (N1802, N1787, N348, N1242, N396);
nor NOR3 (N1803, N1801, N1095, N731);
buf BUF1 (N1804, N1798);
not NOT1 (N1805, N1786);
not NOT1 (N1806, N1803);
and AND2 (N1807, N1783, N348);
and AND4 (N1808, N1804, N1368, N1390, N115);
buf BUF1 (N1809, N1806);
nand NAND2 (N1810, N1800, N1212);
or OR3 (N1811, N1805, N437, N1021);
and AND3 (N1812, N1802, N371, N1050);
and AND2 (N1813, N1808, N260);
buf BUF1 (N1814, N1799);
and AND4 (N1815, N1810, N579, N57, N967);
not NOT1 (N1816, N1807);
xor XOR2 (N1817, N1816, N1496);
not NOT1 (N1818, N1788);
xor XOR2 (N1819, N1813, N208);
not NOT1 (N1820, N1819);
nand NAND2 (N1821, N1817, N1205);
not NOT1 (N1822, N1821);
nand NAND2 (N1823, N1796, N1005);
nor NOR2 (N1824, N1818, N496);
or OR3 (N1825, N1824, N1216, N758);
or OR2 (N1826, N1811, N1512);
nand NAND4 (N1827, N1826, N692, N1178, N184);
buf BUF1 (N1828, N1823);
and AND2 (N1829, N1809, N1713);
nor NOR3 (N1830, N1828, N840, N902);
nand NAND2 (N1831, N1815, N187);
and AND3 (N1832, N1827, N1023, N505);
xor XOR2 (N1833, N1831, N232);
nor NOR2 (N1834, N1832, N1376);
nand NAND2 (N1835, N1825, N685);
and AND4 (N1836, N1820, N745, N1541, N619);
nand NAND2 (N1837, N1829, N161);
xor XOR2 (N1838, N1836, N1454);
and AND4 (N1839, N1834, N334, N940, N1560);
nand NAND2 (N1840, N1822, N314);
and AND3 (N1841, N1812, N686, N1225);
nor NOR2 (N1842, N1814, N1253);
nor NOR4 (N1843, N1797, N1206, N1290, N1793);
xor XOR2 (N1844, N1830, N1284);
nor NOR4 (N1845, N1843, N1768, N469, N73);
xor XOR2 (N1846, N1844, N1703);
nor NOR4 (N1847, N1833, N1519, N87, N244);
and AND2 (N1848, N1838, N1845);
nand NAND2 (N1849, N1496, N83);
or OR3 (N1850, N1835, N1002, N1589);
not NOT1 (N1851, N1850);
xor XOR2 (N1852, N1851, N1428);
not NOT1 (N1853, N1841);
not NOT1 (N1854, N1840);
and AND3 (N1855, N1848, N1112, N1258);
or OR3 (N1856, N1842, N1778, N1577);
and AND2 (N1857, N1853, N1253);
buf BUF1 (N1858, N1854);
and AND4 (N1859, N1858, N764, N1560, N1020);
not NOT1 (N1860, N1852);
nand NAND4 (N1861, N1837, N968, N1419, N719);
and AND4 (N1862, N1847, N1385, N1179, N1557);
nor NOR3 (N1863, N1856, N616, N1384);
and AND2 (N1864, N1846, N402);
nor NOR2 (N1865, N1855, N495);
nor NOR2 (N1866, N1863, N149);
xor XOR2 (N1867, N1862, N1118);
nor NOR3 (N1868, N1839, N1601, N190);
buf BUF1 (N1869, N1866);
buf BUF1 (N1870, N1864);
xor XOR2 (N1871, N1867, N1189);
nand NAND3 (N1872, N1857, N225, N1450);
xor XOR2 (N1873, N1860, N1542);
not NOT1 (N1874, N1868);
not NOT1 (N1875, N1871);
nand NAND2 (N1876, N1875, N1755);
and AND4 (N1877, N1874, N1494, N1767, N1412);
buf BUF1 (N1878, N1873);
xor XOR2 (N1879, N1870, N143);
nor NOR4 (N1880, N1877, N210, N669, N49);
or OR3 (N1881, N1879, N1699, N1151);
nor NOR2 (N1882, N1865, N518);
not NOT1 (N1883, N1859);
and AND2 (N1884, N1861, N1690);
or OR4 (N1885, N1869, N339, N766, N437);
buf BUF1 (N1886, N1882);
or OR2 (N1887, N1886, N691);
and AND4 (N1888, N1880, N351, N942, N765);
xor XOR2 (N1889, N1876, N498);
not NOT1 (N1890, N1881);
and AND2 (N1891, N1849, N852);
nand NAND2 (N1892, N1890, N739);
not NOT1 (N1893, N1872);
nor NOR3 (N1894, N1885, N1582, N726);
nor NOR2 (N1895, N1888, N795);
nand NAND2 (N1896, N1895, N519);
xor XOR2 (N1897, N1887, N1391);
or OR4 (N1898, N1892, N749, N87, N114);
or OR3 (N1899, N1883, N1264, N1526);
or OR2 (N1900, N1893, N746);
not NOT1 (N1901, N1896);
not NOT1 (N1902, N1878);
nor NOR4 (N1903, N1898, N627, N912, N1281);
not NOT1 (N1904, N1902);
xor XOR2 (N1905, N1903, N1877);
not NOT1 (N1906, N1897);
and AND3 (N1907, N1889, N538, N811);
buf BUF1 (N1908, N1907);
or OR3 (N1909, N1905, N718, N1638);
not NOT1 (N1910, N1884);
not NOT1 (N1911, N1900);
or OR3 (N1912, N1904, N410, N1593);
and AND4 (N1913, N1908, N890, N490, N1449);
not NOT1 (N1914, N1910);
buf BUF1 (N1915, N1901);
nor NOR3 (N1916, N1899, N1815, N1412);
not NOT1 (N1917, N1911);
buf BUF1 (N1918, N1912);
buf BUF1 (N1919, N1914);
nand NAND2 (N1920, N1894, N1665);
or OR2 (N1921, N1916, N532);
nand NAND4 (N1922, N1915, N235, N1079, N1359);
nor NOR3 (N1923, N1913, N766, N1336);
nand NAND2 (N1924, N1917, N1163);
not NOT1 (N1925, N1924);
nand NAND2 (N1926, N1918, N1905);
and AND4 (N1927, N1906, N1727, N512, N1376);
buf BUF1 (N1928, N1926);
nand NAND3 (N1929, N1919, N795, N1487);
not NOT1 (N1930, N1929);
and AND2 (N1931, N1928, N1764);
and AND2 (N1932, N1922, N295);
buf BUF1 (N1933, N1921);
not NOT1 (N1934, N1923);
not NOT1 (N1935, N1891);
nor NOR3 (N1936, N1935, N321, N1562);
buf BUF1 (N1937, N1934);
or OR3 (N1938, N1909, N1745, N1645);
xor XOR2 (N1939, N1937, N897);
xor XOR2 (N1940, N1932, N1666);
and AND2 (N1941, N1930, N1135);
nor NOR4 (N1942, N1938, N1137, N880, N1811);
nor NOR4 (N1943, N1936, N1009, N447, N973);
and AND3 (N1944, N1920, N1235, N666);
and AND3 (N1945, N1925, N1228, N1632);
or OR4 (N1946, N1939, N635, N179, N299);
or OR2 (N1947, N1946, N531);
nand NAND2 (N1948, N1945, N1638);
xor XOR2 (N1949, N1943, N1862);
nand NAND3 (N1950, N1933, N1124, N1612);
nor NOR3 (N1951, N1927, N191, N816);
nor NOR3 (N1952, N1949, N1054, N1484);
nand NAND4 (N1953, N1940, N1121, N1236, N1585);
or OR2 (N1954, N1948, N754);
not NOT1 (N1955, N1942);
and AND3 (N1956, N1951, N191, N1164);
xor XOR2 (N1957, N1954, N1149);
nor NOR2 (N1958, N1952, N1156);
xor XOR2 (N1959, N1947, N847);
buf BUF1 (N1960, N1958);
or OR2 (N1961, N1959, N1637);
xor XOR2 (N1962, N1950, N209);
nor NOR3 (N1963, N1960, N34, N310);
nor NOR2 (N1964, N1957, N623);
buf BUF1 (N1965, N1962);
and AND2 (N1966, N1941, N1929);
xor XOR2 (N1967, N1964, N1546);
buf BUF1 (N1968, N1965);
xor XOR2 (N1969, N1968, N1848);
not NOT1 (N1970, N1961);
not NOT1 (N1971, N1956);
not NOT1 (N1972, N1963);
nor NOR4 (N1973, N1944, N259, N1244, N1730);
nor NOR2 (N1974, N1972, N564);
buf BUF1 (N1975, N1969);
nand NAND4 (N1976, N1974, N609, N388, N817);
and AND4 (N1977, N1975, N1566, N1327, N1889);
buf BUF1 (N1978, N1966);
not NOT1 (N1979, N1955);
nor NOR3 (N1980, N1970, N1255, N1198);
buf BUF1 (N1981, N1973);
not NOT1 (N1982, N1981);
nor NOR3 (N1983, N1979, N1821, N601);
nor NOR2 (N1984, N1978, N727);
and AND3 (N1985, N1971, N1381, N334);
or OR4 (N1986, N1984, N775, N1240, N337);
nand NAND4 (N1987, N1931, N1108, N415, N757);
nand NAND4 (N1988, N1976, N620, N500, N1558);
and AND4 (N1989, N1986, N1929, N1570, N252);
not NOT1 (N1990, N1977);
nor NOR3 (N1991, N1988, N674, N880);
nand NAND2 (N1992, N1991, N1718);
and AND2 (N1993, N1982, N1606);
and AND4 (N1994, N1980, N976, N247, N198);
nor NOR4 (N1995, N1993, N1585, N167, N1624);
nor NOR4 (N1996, N1983, N253, N429, N787);
or OR4 (N1997, N1987, N1928, N849, N376);
not NOT1 (N1998, N1990);
not NOT1 (N1999, N1989);
buf BUF1 (N2000, N1997);
xor XOR2 (N2001, N1999, N1352);
not NOT1 (N2002, N1998);
nand NAND2 (N2003, N2002, N854);
nand NAND3 (N2004, N1994, N1455, N964);
buf BUF1 (N2005, N2001);
buf BUF1 (N2006, N1953);
nand NAND3 (N2007, N1992, N1003, N1957);
nor NOR4 (N2008, N2006, N1377, N722, N397);
xor XOR2 (N2009, N1967, N1388);
xor XOR2 (N2010, N2000, N20);
and AND4 (N2011, N1985, N8, N1882, N1012);
buf BUF1 (N2012, N2007);
buf BUF1 (N2013, N2003);
buf BUF1 (N2014, N2011);
and AND3 (N2015, N2005, N1145, N1539);
xor XOR2 (N2016, N1995, N473);
and AND4 (N2017, N2008, N1920, N1141, N151);
and AND4 (N2018, N2014, N1269, N1718, N1512);
nor NOR2 (N2019, N2018, N1032);
and AND3 (N2020, N2010, N539, N90);
and AND2 (N2021, N2016, N1663);
not NOT1 (N2022, N2021);
and AND2 (N2023, N2019, N1381);
xor XOR2 (N2024, N1996, N2004);
buf BUF1 (N2025, N444);
or OR2 (N2026, N2009, N340);
buf BUF1 (N2027, N2024);
nand NAND4 (N2028, N2012, N1347, N1634, N1523);
xor XOR2 (N2029, N2026, N1543);
and AND4 (N2030, N2022, N1021, N1552, N506);
nand NAND3 (N2031, N2029, N297, N422);
or OR3 (N2032, N2013, N609, N999);
xor XOR2 (N2033, N2025, N661);
not NOT1 (N2034, N2020);
nor NOR3 (N2035, N2015, N773, N1418);
xor XOR2 (N2036, N2033, N892);
or OR3 (N2037, N2034, N1721, N418);
buf BUF1 (N2038, N2037);
buf BUF1 (N2039, N2030);
xor XOR2 (N2040, N2032, N1425);
nor NOR4 (N2041, N2028, N1245, N1839, N1993);
nor NOR3 (N2042, N2031, N1298, N1801);
nand NAND4 (N2043, N2039, N78, N333, N733);
nor NOR3 (N2044, N2036, N1325, N1833);
and AND4 (N2045, N2040, N1568, N190, N1783);
not NOT1 (N2046, N2035);
nor NOR3 (N2047, N2045, N407, N222);
and AND4 (N2048, N2023, N287, N1404, N1561);
and AND3 (N2049, N2043, N1358, N1321);
buf BUF1 (N2050, N2027);
nand NAND3 (N2051, N2038, N1459, N1262);
not NOT1 (N2052, N2017);
xor XOR2 (N2053, N2044, N350);
xor XOR2 (N2054, N2041, N1684);
nand NAND3 (N2055, N2042, N320, N341);
not NOT1 (N2056, N2050);
nand NAND2 (N2057, N2049, N553);
and AND4 (N2058, N2056, N1222, N311, N1830);
nand NAND2 (N2059, N2051, N1075);
not NOT1 (N2060, N2047);
xor XOR2 (N2061, N2052, N2045);
and AND2 (N2062, N2046, N1305);
xor XOR2 (N2063, N2057, N1057);
and AND2 (N2064, N2059, N1633);
nor NOR3 (N2065, N2053, N986, N1843);
and AND2 (N2066, N2048, N1940);
or OR3 (N2067, N2060, N1192, N2055);
or OR2 (N2068, N1919, N1987);
nor NOR2 (N2069, N2066, N160);
nand NAND2 (N2070, N2063, N289);
and AND2 (N2071, N2062, N1269);
or OR3 (N2072, N2064, N703, N480);
and AND3 (N2073, N2054, N1268, N417);
nor NOR3 (N2074, N2068, N849, N1234);
and AND3 (N2075, N2065, N825, N1869);
xor XOR2 (N2076, N2067, N770);
buf BUF1 (N2077, N2070);
or OR3 (N2078, N2058, N1270, N1174);
buf BUF1 (N2079, N2069);
nand NAND4 (N2080, N2061, N178, N720, N1589);
not NOT1 (N2081, N2076);
xor XOR2 (N2082, N2075, N52);
or OR4 (N2083, N2071, N147, N1154, N730);
xor XOR2 (N2084, N2082, N1451);
and AND2 (N2085, N2078, N1195);
buf BUF1 (N2086, N2073);
and AND3 (N2087, N2081, N262, N2083);
not NOT1 (N2088, N968);
or OR4 (N2089, N2074, N1077, N1799, N1084);
buf BUF1 (N2090, N2077);
nor NOR4 (N2091, N2080, N1255, N1996, N1175);
or OR3 (N2092, N2072, N1306, N1500);
xor XOR2 (N2093, N2088, N751);
or OR3 (N2094, N2092, N84, N879);
nand NAND3 (N2095, N2089, N2015, N890);
xor XOR2 (N2096, N2087, N505);
and AND2 (N2097, N2084, N1234);
buf BUF1 (N2098, N2095);
nor NOR2 (N2099, N2086, N1391);
xor XOR2 (N2100, N2097, N259);
nand NAND3 (N2101, N2093, N1275, N1822);
nor NOR2 (N2102, N2091, N1894);
nand NAND2 (N2103, N2090, N1151);
and AND4 (N2104, N2094, N648, N487, N193);
nand NAND3 (N2105, N2100, N850, N515);
nand NAND3 (N2106, N2079, N482, N1222);
and AND4 (N2107, N2106, N1971, N143, N475);
not NOT1 (N2108, N2085);
and AND2 (N2109, N2099, N1814);
nor NOR4 (N2110, N2104, N722, N226, N2062);
and AND2 (N2111, N2105, N730);
or OR3 (N2112, N2110, N672, N829);
not NOT1 (N2113, N2096);
and AND3 (N2114, N2107, N788, N31);
nand NAND3 (N2115, N2113, N1001, N1999);
xor XOR2 (N2116, N2114, N63);
nand NAND3 (N2117, N2111, N1261, N835);
or OR4 (N2118, N2108, N242, N834, N264);
or OR3 (N2119, N2098, N1180, N1880);
nor NOR4 (N2120, N2102, N862, N721, N1321);
nand NAND2 (N2121, N2109, N347);
xor XOR2 (N2122, N2115, N104);
or OR4 (N2123, N2116, N1415, N1091, N1241);
buf BUF1 (N2124, N2118);
nand NAND2 (N2125, N2123, N510);
buf BUF1 (N2126, N2121);
and AND3 (N2127, N2101, N1787, N937);
and AND2 (N2128, N2112, N61);
xor XOR2 (N2129, N2125, N1523);
or OR3 (N2130, N2126, N651, N32);
or OR4 (N2131, N2124, N771, N175, N425);
or OR2 (N2132, N2131, N764);
xor XOR2 (N2133, N2120, N1782);
xor XOR2 (N2134, N2133, N694);
not NOT1 (N2135, N2134);
and AND4 (N2136, N2132, N1442, N1411, N1846);
not NOT1 (N2137, N2135);
nor NOR4 (N2138, N2129, N830, N872, N1065);
buf BUF1 (N2139, N2138);
xor XOR2 (N2140, N2139, N803);
buf BUF1 (N2141, N2119);
not NOT1 (N2142, N2122);
buf BUF1 (N2143, N2130);
nand NAND2 (N2144, N2103, N1276);
nor NOR4 (N2145, N2136, N620, N450, N1395);
not NOT1 (N2146, N2127);
and AND3 (N2147, N2143, N1458, N118);
xor XOR2 (N2148, N2144, N1670);
xor XOR2 (N2149, N2142, N1490);
nand NAND4 (N2150, N2117, N1358, N620, N346);
buf BUF1 (N2151, N2141);
buf BUF1 (N2152, N2128);
nand NAND2 (N2153, N2152, N998);
and AND2 (N2154, N2151, N1821);
buf BUF1 (N2155, N2148);
nor NOR2 (N2156, N2155, N653);
nor NOR2 (N2157, N2140, N7);
and AND2 (N2158, N2150, N690);
not NOT1 (N2159, N2154);
nor NOR4 (N2160, N2147, N1623, N2111, N155);
or OR3 (N2161, N2145, N3, N879);
and AND4 (N2162, N2159, N2025, N861, N1938);
not NOT1 (N2163, N2156);
buf BUF1 (N2164, N2163);
xor XOR2 (N2165, N2146, N1727);
or OR4 (N2166, N2137, N21, N781, N1007);
buf BUF1 (N2167, N2160);
nor NOR4 (N2168, N2158, N1162, N2146, N868);
buf BUF1 (N2169, N2167);
nor NOR3 (N2170, N2165, N816, N1229);
not NOT1 (N2171, N2169);
and AND3 (N2172, N2164, N250, N1035);
xor XOR2 (N2173, N2166, N1249);
or OR3 (N2174, N2162, N1842, N2159);
xor XOR2 (N2175, N2171, N1618);
buf BUF1 (N2176, N2172);
and AND2 (N2177, N2173, N619);
nand NAND3 (N2178, N2157, N834, N1594);
xor XOR2 (N2179, N2176, N446);
or OR4 (N2180, N2178, N1317, N1800, N2032);
or OR2 (N2181, N2149, N1246);
buf BUF1 (N2182, N2170);
xor XOR2 (N2183, N2181, N454);
xor XOR2 (N2184, N2153, N1512);
nor NOR4 (N2185, N2174, N106, N1774, N1792);
nand NAND2 (N2186, N2179, N1325);
or OR2 (N2187, N2186, N1227);
xor XOR2 (N2188, N2180, N1326);
and AND3 (N2189, N2187, N607, N1146);
and AND4 (N2190, N2175, N1929, N1662, N2182);
nor NOR3 (N2191, N16, N522, N48);
not NOT1 (N2192, N2185);
buf BUF1 (N2193, N2184);
nand NAND2 (N2194, N2183, N2143);
buf BUF1 (N2195, N2193);
or OR3 (N2196, N2188, N1364, N1582);
xor XOR2 (N2197, N2192, N1369);
nor NOR2 (N2198, N2189, N47);
xor XOR2 (N2199, N2168, N1005);
nand NAND2 (N2200, N2195, N1215);
and AND2 (N2201, N2200, N91);
nor NOR2 (N2202, N2198, N2037);
not NOT1 (N2203, N2161);
xor XOR2 (N2204, N2197, N1293);
buf BUF1 (N2205, N2201);
nor NOR4 (N2206, N2191, N2153, N901, N1552);
not NOT1 (N2207, N2194);
not NOT1 (N2208, N2196);
not NOT1 (N2209, N2199);
and AND3 (N2210, N2204, N205, N2066);
and AND4 (N2211, N2209, N296, N274, N1285);
nand NAND2 (N2212, N2210, N110);
buf BUF1 (N2213, N2211);
buf BUF1 (N2214, N2213);
and AND2 (N2215, N2208, N723);
not NOT1 (N2216, N2190);
buf BUF1 (N2217, N2206);
buf BUF1 (N2218, N2202);
and AND3 (N2219, N2203, N1855, N942);
nand NAND3 (N2220, N2205, N412, N1984);
buf BUF1 (N2221, N2216);
and AND4 (N2222, N2217, N470, N1886, N1784);
nor NOR4 (N2223, N2220, N913, N2164, N626);
and AND2 (N2224, N2219, N821);
nor NOR3 (N2225, N2212, N693, N412);
not NOT1 (N2226, N2214);
and AND3 (N2227, N2225, N786, N1314);
not NOT1 (N2228, N2222);
or OR3 (N2229, N2215, N364, N1190);
nor NOR4 (N2230, N2207, N476, N1323, N1079);
not NOT1 (N2231, N2229);
and AND3 (N2232, N2231, N545, N2227);
or OR4 (N2233, N1081, N251, N655, N506);
or OR4 (N2234, N2232, N1661, N59, N2100);
nor NOR3 (N2235, N2224, N1209, N1153);
or OR4 (N2236, N2226, N1846, N899, N1298);
buf BUF1 (N2237, N2223);
buf BUF1 (N2238, N2218);
and AND3 (N2239, N2221, N724, N1005);
nor NOR4 (N2240, N2234, N246, N762, N1034);
xor XOR2 (N2241, N2235, N437);
xor XOR2 (N2242, N2238, N1416);
or OR3 (N2243, N2242, N529, N1672);
buf BUF1 (N2244, N2239);
nor NOR2 (N2245, N2244, N1120);
nand NAND3 (N2246, N2233, N267, N1306);
buf BUF1 (N2247, N2236);
and AND3 (N2248, N2245, N1835, N1108);
not NOT1 (N2249, N2230);
xor XOR2 (N2250, N2241, N148);
or OR2 (N2251, N2248, N2175);
or OR3 (N2252, N2228, N114, N561);
not NOT1 (N2253, N2240);
nand NAND3 (N2254, N2250, N361, N1029);
nand NAND3 (N2255, N2177, N384, N1552);
or OR3 (N2256, N2246, N3, N1040);
and AND2 (N2257, N2249, N1147);
and AND4 (N2258, N2243, N1184, N2163, N1186);
nor NOR3 (N2259, N2255, N1652, N1961);
nor NOR3 (N2260, N2247, N781, N137);
not NOT1 (N2261, N2253);
nand NAND2 (N2262, N2256, N738);
xor XOR2 (N2263, N2258, N2045);
and AND2 (N2264, N2254, N1281);
and AND4 (N2265, N2264, N1266, N1784, N365);
and AND2 (N2266, N2262, N173);
nand NAND2 (N2267, N2257, N790);
nand NAND3 (N2268, N2260, N2078, N1187);
nor NOR4 (N2269, N2267, N729, N2226, N1049);
and AND4 (N2270, N2269, N1875, N2149, N2221);
buf BUF1 (N2271, N2261);
or OR3 (N2272, N2263, N92, N1619);
not NOT1 (N2273, N2251);
and AND3 (N2274, N2273, N628, N2086);
nand NAND3 (N2275, N2270, N1093, N971);
not NOT1 (N2276, N2265);
and AND3 (N2277, N2272, N578, N914);
not NOT1 (N2278, N2274);
nand NAND2 (N2279, N2268, N1533);
xor XOR2 (N2280, N2276, N790);
not NOT1 (N2281, N2259);
or OR4 (N2282, N2275, N115, N1445, N323);
and AND2 (N2283, N2252, N882);
buf BUF1 (N2284, N2282);
not NOT1 (N2285, N2277);
xor XOR2 (N2286, N2266, N639);
not NOT1 (N2287, N2286);
buf BUF1 (N2288, N2237);
nand NAND2 (N2289, N2278, N1335);
xor XOR2 (N2290, N2285, N1061);
xor XOR2 (N2291, N2281, N1710);
buf BUF1 (N2292, N2284);
xor XOR2 (N2293, N2292, N1227);
not NOT1 (N2294, N2288);
buf BUF1 (N2295, N2279);
nor NOR4 (N2296, N2289, N1758, N1929, N877);
or OR2 (N2297, N2293, N763);
nor NOR4 (N2298, N2295, N2229, N849, N1285);
buf BUF1 (N2299, N2283);
not NOT1 (N2300, N2291);
or OR2 (N2301, N2271, N1222);
nand NAND4 (N2302, N2287, N237, N548, N48);
nor NOR3 (N2303, N2297, N1578, N1090);
and AND2 (N2304, N2298, N861);
or OR4 (N2305, N2300, N1642, N29, N471);
or OR4 (N2306, N2304, N1220, N1459, N985);
and AND3 (N2307, N2305, N1717, N1612);
xor XOR2 (N2308, N2307, N1171);
xor XOR2 (N2309, N2280, N1651);
or OR3 (N2310, N2294, N1452, N502);
xor XOR2 (N2311, N2299, N1836);
not NOT1 (N2312, N2308);
or OR3 (N2313, N2306, N833, N79);
xor XOR2 (N2314, N2296, N1832);
xor XOR2 (N2315, N2311, N1475);
and AND4 (N2316, N2314, N1312, N785, N672);
xor XOR2 (N2317, N2310, N227);
xor XOR2 (N2318, N2313, N650);
nor NOR4 (N2319, N2315, N1496, N929, N659);
nor NOR4 (N2320, N2317, N576, N2166, N746);
and AND2 (N2321, N2312, N69);
xor XOR2 (N2322, N2302, N1480);
nor NOR3 (N2323, N2319, N1454, N47);
nand NAND3 (N2324, N2303, N1695, N1997);
nand NAND4 (N2325, N2324, N2203, N1155, N1113);
and AND2 (N2326, N2322, N2156);
or OR4 (N2327, N2321, N1967, N1268, N1070);
buf BUF1 (N2328, N2318);
nand NAND2 (N2329, N2316, N387);
or OR3 (N2330, N2327, N1382, N1349);
xor XOR2 (N2331, N2323, N1326);
xor XOR2 (N2332, N2325, N1860);
or OR4 (N2333, N2290, N481, N330, N279);
nand NAND3 (N2334, N2309, N1561, N313);
xor XOR2 (N2335, N2332, N1467);
and AND2 (N2336, N2331, N448);
or OR2 (N2337, N2326, N1869);
not NOT1 (N2338, N2334);
or OR4 (N2339, N2330, N839, N136, N563);
not NOT1 (N2340, N2333);
nand NAND4 (N2341, N2336, N961, N2084, N851);
and AND2 (N2342, N2328, N1510);
or OR4 (N2343, N2341, N508, N2187, N1250);
or OR2 (N2344, N2338, N2245);
or OR3 (N2345, N2344, N853, N225);
nor NOR3 (N2346, N2340, N1279, N1749);
nor NOR3 (N2347, N2339, N316, N1297);
nand NAND4 (N2348, N2337, N1763, N2192, N1407);
nor NOR2 (N2349, N2342, N797);
and AND4 (N2350, N2345, N2329, N317, N361);
not NOT1 (N2351, N292);
not NOT1 (N2352, N2343);
and AND2 (N2353, N2350, N450);
nor NOR4 (N2354, N2348, N594, N1562, N1638);
nand NAND4 (N2355, N2346, N85, N132, N830);
xor XOR2 (N2356, N2320, N1756);
nor NOR3 (N2357, N2301, N570, N999);
nand NAND4 (N2358, N2352, N132, N385, N1061);
buf BUF1 (N2359, N2354);
or OR4 (N2360, N2349, N992, N432, N1008);
nand NAND3 (N2361, N2353, N393, N1315);
buf BUF1 (N2362, N2355);
xor XOR2 (N2363, N2335, N1080);
not NOT1 (N2364, N2362);
nand NAND2 (N2365, N2347, N2113);
not NOT1 (N2366, N2363);
or OR4 (N2367, N2359, N393, N335, N541);
not NOT1 (N2368, N2351);
xor XOR2 (N2369, N2366, N115);
xor XOR2 (N2370, N2368, N1420);
nand NAND4 (N2371, N2370, N1344, N1808, N2292);
nor NOR2 (N2372, N2356, N22);
nand NAND3 (N2373, N2367, N1225, N252);
buf BUF1 (N2374, N2371);
nand NAND4 (N2375, N2372, N246, N1747, N109);
or OR2 (N2376, N2375, N1390);
not NOT1 (N2377, N2369);
xor XOR2 (N2378, N2373, N2085);
and AND2 (N2379, N2361, N583);
not NOT1 (N2380, N2365);
nor NOR2 (N2381, N2379, N1380);
xor XOR2 (N2382, N2380, N1666);
not NOT1 (N2383, N2357);
and AND4 (N2384, N2378, N1105, N516, N366);
and AND4 (N2385, N2358, N614, N1534, N600);
nand NAND3 (N2386, N2364, N312, N967);
not NOT1 (N2387, N2377);
not NOT1 (N2388, N2386);
xor XOR2 (N2389, N2388, N1476);
nand NAND2 (N2390, N2360, N43);
and AND3 (N2391, N2374, N1717, N275);
not NOT1 (N2392, N2385);
buf BUF1 (N2393, N2391);
nor NOR2 (N2394, N2384, N505);
not NOT1 (N2395, N2389);
or OR2 (N2396, N2390, N174);
and AND2 (N2397, N2394, N342);
nor NOR4 (N2398, N2376, N1104, N1490, N1496);
nand NAND3 (N2399, N2382, N1822, N962);
and AND2 (N2400, N2381, N614);
xor XOR2 (N2401, N2396, N935);
nand NAND4 (N2402, N2395, N519, N679, N1438);
buf BUF1 (N2403, N2401);
and AND4 (N2404, N2392, N405, N1335, N419);
buf BUF1 (N2405, N2400);
nand NAND3 (N2406, N2383, N1285, N737);
or OR2 (N2407, N2387, N2086);
nor NOR2 (N2408, N2397, N829);
xor XOR2 (N2409, N2405, N263);
nand NAND2 (N2410, N2399, N923);
buf BUF1 (N2411, N2407);
buf BUF1 (N2412, N2404);
buf BUF1 (N2413, N2406);
buf BUF1 (N2414, N2409);
or OR4 (N2415, N2413, N854, N870, N520);
xor XOR2 (N2416, N2398, N1732);
not NOT1 (N2417, N2415);
nor NOR4 (N2418, N2411, N2385, N515, N1060);
nand NAND2 (N2419, N2417, N1556);
xor XOR2 (N2420, N2418, N180);
or OR3 (N2421, N2402, N394, N171);
xor XOR2 (N2422, N2410, N1514);
xor XOR2 (N2423, N2393, N657);
nor NOR2 (N2424, N2414, N1294);
xor XOR2 (N2425, N2421, N179);
nor NOR4 (N2426, N2408, N2252, N1370, N2193);
not NOT1 (N2427, N2423);
buf BUF1 (N2428, N2412);
buf BUF1 (N2429, N2425);
nand NAND2 (N2430, N2419, N2061);
xor XOR2 (N2431, N2424, N214);
xor XOR2 (N2432, N2428, N1429);
buf BUF1 (N2433, N2427);
buf BUF1 (N2434, N2426);
or OR4 (N2435, N2431, N1047, N1832, N1239);
buf BUF1 (N2436, N2420);
nor NOR3 (N2437, N2435, N1044, N235);
or OR4 (N2438, N2432, N1419, N1725, N1769);
and AND4 (N2439, N2433, N242, N2423, N2419);
buf BUF1 (N2440, N2434);
or OR4 (N2441, N2422, N2322, N1130, N350);
nand NAND3 (N2442, N2437, N573, N1914);
and AND3 (N2443, N2442, N1702, N1577);
xor XOR2 (N2444, N2403, N2384);
xor XOR2 (N2445, N2440, N2064);
not NOT1 (N2446, N2444);
not NOT1 (N2447, N2438);
xor XOR2 (N2448, N2445, N176);
not NOT1 (N2449, N2448);
buf BUF1 (N2450, N2430);
nand NAND2 (N2451, N2441, N1046);
nand NAND3 (N2452, N2439, N1199, N1608);
nand NAND4 (N2453, N2446, N1546, N1783, N1017);
nor NOR3 (N2454, N2452, N1437, N587);
and AND3 (N2455, N2450, N1765, N1418);
buf BUF1 (N2456, N2455);
nand NAND3 (N2457, N2449, N964, N1347);
nor NOR2 (N2458, N2443, N870);
buf BUF1 (N2459, N2451);
nor NOR3 (N2460, N2447, N2429, N1120);
not NOT1 (N2461, N604);
nor NOR4 (N2462, N2460, N914, N819, N2163);
and AND3 (N2463, N2457, N1671, N706);
or OR3 (N2464, N2462, N2456, N1319);
xor XOR2 (N2465, N333, N1161);
and AND2 (N2466, N2461, N378);
or OR3 (N2467, N2458, N1018, N2428);
and AND2 (N2468, N2463, N2043);
xor XOR2 (N2469, N2466, N1191);
nand NAND2 (N2470, N2453, N1006);
nor NOR2 (N2471, N2465, N2437);
xor XOR2 (N2472, N2459, N1337);
xor XOR2 (N2473, N2464, N1209);
nor NOR2 (N2474, N2470, N779);
buf BUF1 (N2475, N2469);
nand NAND2 (N2476, N2472, N433);
nor NOR3 (N2477, N2473, N1350, N1981);
xor XOR2 (N2478, N2454, N286);
or OR2 (N2479, N2416, N728);
nor NOR4 (N2480, N2475, N741, N34, N1314);
not NOT1 (N2481, N2476);
nor NOR2 (N2482, N2467, N1599);
buf BUF1 (N2483, N2481);
xor XOR2 (N2484, N2478, N471);
nor NOR2 (N2485, N2482, N329);
or OR4 (N2486, N2483, N273, N1008, N1149);
buf BUF1 (N2487, N2436);
nand NAND2 (N2488, N2487, N224);
buf BUF1 (N2489, N2474);
nor NOR4 (N2490, N2477, N675, N23, N2251);
and AND2 (N2491, N2490, N1066);
not NOT1 (N2492, N2486);
nor NOR4 (N2493, N2468, N2366, N337, N2322);
or OR3 (N2494, N2489, N813, N685);
and AND2 (N2495, N2488, N1913);
or OR4 (N2496, N2485, N1954, N1441, N654);
nor NOR4 (N2497, N2491, N1991, N1377, N791);
and AND2 (N2498, N2492, N706);
or OR4 (N2499, N2471, N105, N1970, N1455);
or OR3 (N2500, N2497, N1772, N2299);
and AND4 (N2501, N2484, N512, N1739, N431);
or OR3 (N2502, N2493, N2117, N996);
and AND3 (N2503, N2479, N2271, N326);
and AND4 (N2504, N2503, N1884, N2396, N1293);
not NOT1 (N2505, N2500);
not NOT1 (N2506, N2501);
nand NAND3 (N2507, N2498, N1182, N656);
or OR4 (N2508, N2507, N1257, N1165, N2232);
and AND2 (N2509, N2504, N887);
buf BUF1 (N2510, N2508);
buf BUF1 (N2511, N2499);
nor NOR3 (N2512, N2480, N794, N526);
nand NAND3 (N2513, N2502, N100, N514);
buf BUF1 (N2514, N2509);
or OR3 (N2515, N2511, N1222, N102);
or OR3 (N2516, N2512, N1935, N2160);
not NOT1 (N2517, N2496);
buf BUF1 (N2518, N2517);
buf BUF1 (N2519, N2516);
and AND2 (N2520, N2506, N577);
or OR2 (N2521, N2514, N1488);
or OR3 (N2522, N2521, N292, N1854);
or OR3 (N2523, N2522, N2370, N730);
xor XOR2 (N2524, N2523, N284);
nand NAND4 (N2525, N2494, N245, N2323, N839);
or OR3 (N2526, N2524, N1487, N2485);
nand NAND2 (N2527, N2519, N2352);
nor NOR2 (N2528, N2515, N2);
and AND2 (N2529, N2525, N1891);
or OR3 (N2530, N2527, N1758, N1877);
nand NAND4 (N2531, N2530, N945, N1751, N1957);
buf BUF1 (N2532, N2513);
nor NOR2 (N2533, N2510, N1066);
and AND4 (N2534, N2495, N281, N1177, N487);
or OR4 (N2535, N2528, N296, N1108, N1216);
nor NOR4 (N2536, N2532, N1996, N1878, N563);
xor XOR2 (N2537, N2535, N261);
or OR2 (N2538, N2505, N190);
and AND4 (N2539, N2526, N1269, N2045, N1678);
and AND3 (N2540, N2536, N2288, N692);
buf BUF1 (N2541, N2540);
buf BUF1 (N2542, N2533);
nor NOR4 (N2543, N2520, N1160, N1694, N1056);
xor XOR2 (N2544, N2538, N920);
xor XOR2 (N2545, N2529, N2320);
and AND2 (N2546, N2545, N2090);
nor NOR2 (N2547, N2541, N746);
xor XOR2 (N2548, N2547, N1335);
and AND2 (N2549, N2518, N1063);
nor NOR4 (N2550, N2548, N1514, N2321, N2023);
nor NOR3 (N2551, N2550, N580, N849);
not NOT1 (N2552, N2531);
not NOT1 (N2553, N2546);
and AND4 (N2554, N2537, N990, N1242, N2313);
nor NOR4 (N2555, N2544, N2267, N2500, N1489);
xor XOR2 (N2556, N2551, N2030);
nand NAND4 (N2557, N2555, N1020, N1237, N1863);
nand NAND3 (N2558, N2543, N779, N2306);
and AND3 (N2559, N2554, N793, N2527);
xor XOR2 (N2560, N2534, N766);
and AND2 (N2561, N2558, N1242);
and AND3 (N2562, N2560, N2512, N1188);
xor XOR2 (N2563, N2556, N1091);
xor XOR2 (N2564, N2559, N1545);
xor XOR2 (N2565, N2561, N1629);
and AND4 (N2566, N2557, N748, N1303, N1783);
and AND4 (N2567, N2539, N347, N290, N2041);
xor XOR2 (N2568, N2564, N1642);
or OR2 (N2569, N2562, N172);
and AND3 (N2570, N2549, N167, N2527);
xor XOR2 (N2571, N2553, N750);
or OR4 (N2572, N2569, N859, N1069, N759);
buf BUF1 (N2573, N2552);
buf BUF1 (N2574, N2563);
not NOT1 (N2575, N2567);
nand NAND4 (N2576, N2572, N625, N1057, N1865);
and AND2 (N2577, N2566, N186);
not NOT1 (N2578, N2575);
not NOT1 (N2579, N2573);
nor NOR2 (N2580, N2579, N572);
or OR4 (N2581, N2542, N1535, N1922, N202);
xor XOR2 (N2582, N2570, N828);
not NOT1 (N2583, N2577);
nor NOR3 (N2584, N2565, N1749, N1798);
not NOT1 (N2585, N2576);
nand NAND2 (N2586, N2582, N982);
buf BUF1 (N2587, N2574);
nand NAND2 (N2588, N2586, N1100);
not NOT1 (N2589, N2583);
nand NAND3 (N2590, N2580, N1995, N1960);
buf BUF1 (N2591, N2578);
nand NAND4 (N2592, N2589, N2082, N150, N465);
not NOT1 (N2593, N2585);
not NOT1 (N2594, N2592);
not NOT1 (N2595, N2584);
xor XOR2 (N2596, N2590, N2477);
and AND4 (N2597, N2591, N1738, N1323, N586);
nand NAND4 (N2598, N2581, N217, N1552, N957);
xor XOR2 (N2599, N2598, N1659);
xor XOR2 (N2600, N2597, N638);
not NOT1 (N2601, N2599);
xor XOR2 (N2602, N2600, N1045);
or OR2 (N2603, N2596, N1912);
nand NAND3 (N2604, N2594, N305, N156);
nand NAND2 (N2605, N2593, N1230);
buf BUF1 (N2606, N2571);
buf BUF1 (N2607, N2603);
nand NAND4 (N2608, N2568, N209, N78, N65);
nor NOR3 (N2609, N2601, N1012, N427);
xor XOR2 (N2610, N2595, N344);
or OR3 (N2611, N2602, N1413, N729);
or OR4 (N2612, N2606, N1196, N1629, N1223);
xor XOR2 (N2613, N2588, N1953);
and AND3 (N2614, N2613, N2437, N183);
nand NAND3 (N2615, N2614, N1381, N2394);
xor XOR2 (N2616, N2608, N2614);
xor XOR2 (N2617, N2609, N816);
nand NAND4 (N2618, N2587, N882, N65, N2309);
or OR4 (N2619, N2607, N1691, N1622, N2311);
buf BUF1 (N2620, N2605);
nor NOR4 (N2621, N2604, N2244, N572, N1378);
and AND3 (N2622, N2612, N867, N892);
buf BUF1 (N2623, N2618);
or OR2 (N2624, N2611, N618);
buf BUF1 (N2625, N2622);
not NOT1 (N2626, N2615);
nand NAND2 (N2627, N2625, N2374);
and AND2 (N2628, N2620, N1601);
xor XOR2 (N2629, N2626, N1358);
xor XOR2 (N2630, N2629, N2461);
nand NAND3 (N2631, N2624, N994, N2314);
not NOT1 (N2632, N2610);
not NOT1 (N2633, N2628);
xor XOR2 (N2634, N2621, N683);
buf BUF1 (N2635, N2634);
not NOT1 (N2636, N2619);
and AND2 (N2637, N2633, N2577);
or OR2 (N2638, N2616, N2300);
or OR3 (N2639, N2630, N952, N1756);
or OR2 (N2640, N2638, N2165);
or OR3 (N2641, N2631, N2424, N63);
xor XOR2 (N2642, N2627, N1776);
nor NOR4 (N2643, N2617, N1082, N2247, N566);
buf BUF1 (N2644, N2623);
xor XOR2 (N2645, N2635, N949);
or OR2 (N2646, N2636, N1025);
not NOT1 (N2647, N2645);
nor NOR4 (N2648, N2639, N377, N1191, N130);
and AND2 (N2649, N2644, N634);
and AND4 (N2650, N2649, N1401, N2531, N1715);
nor NOR3 (N2651, N2643, N1886, N638);
not NOT1 (N2652, N2640);
or OR2 (N2653, N2641, N842);
or OR2 (N2654, N2647, N704);
nand NAND3 (N2655, N2650, N1742, N1460);
not NOT1 (N2656, N2651);
and AND2 (N2657, N2654, N525);
or OR2 (N2658, N2657, N164);
and AND4 (N2659, N2656, N2457, N514, N2629);
buf BUF1 (N2660, N2652);
and AND4 (N2661, N2655, N2588, N1047, N2042);
nor NOR3 (N2662, N2648, N1626, N2313);
buf BUF1 (N2663, N2658);
not NOT1 (N2664, N2646);
not NOT1 (N2665, N2637);
xor XOR2 (N2666, N2632, N2355);
not NOT1 (N2667, N2653);
xor XOR2 (N2668, N2642, N466);
and AND2 (N2669, N2660, N2151);
nand NAND2 (N2670, N2668, N2384);
and AND3 (N2671, N2665, N2153, N1175);
xor XOR2 (N2672, N2667, N809);
nor NOR3 (N2673, N2659, N1503, N1443);
buf BUF1 (N2674, N2663);
and AND3 (N2675, N2666, N451, N36);
or OR3 (N2676, N2664, N2251, N2375);
not NOT1 (N2677, N2676);
not NOT1 (N2678, N2670);
xor XOR2 (N2679, N2678, N2387);
xor XOR2 (N2680, N2679, N782);
nand NAND2 (N2681, N2677, N758);
buf BUF1 (N2682, N2672);
and AND4 (N2683, N2682, N1768, N1739, N2495);
and AND3 (N2684, N2671, N2304, N660);
xor XOR2 (N2685, N2669, N267);
not NOT1 (N2686, N2683);
nand NAND3 (N2687, N2681, N1964, N2407);
buf BUF1 (N2688, N2661);
not NOT1 (N2689, N2680);
or OR2 (N2690, N2673, N454);
xor XOR2 (N2691, N2685, N2350);
nor NOR2 (N2692, N2691, N1255);
nand NAND2 (N2693, N2688, N847);
and AND2 (N2694, N2674, N830);
nand NAND3 (N2695, N2690, N1457, N625);
nor NOR2 (N2696, N2692, N1634);
buf BUF1 (N2697, N2694);
and AND3 (N2698, N2687, N1745, N701);
xor XOR2 (N2699, N2697, N1241);
not NOT1 (N2700, N2684);
buf BUF1 (N2701, N2662);
buf BUF1 (N2702, N2699);
or OR3 (N2703, N2700, N611, N1988);
and AND4 (N2704, N2698, N202, N2017, N1220);
not NOT1 (N2705, N2695);
nor NOR2 (N2706, N2686, N2462);
and AND2 (N2707, N2705, N743);
not NOT1 (N2708, N2675);
nand NAND4 (N2709, N2707, N79, N2396, N1736);
and AND4 (N2710, N2689, N639, N1017, N406);
buf BUF1 (N2711, N2708);
xor XOR2 (N2712, N2693, N40);
and AND3 (N2713, N2701, N1725, N2306);
nor NOR3 (N2714, N2696, N972, N2452);
not NOT1 (N2715, N2714);
buf BUF1 (N2716, N2702);
nand NAND4 (N2717, N2712, N2308, N705, N92);
nor NOR3 (N2718, N2709, N2090, N664);
nor NOR4 (N2719, N2710, N2040, N972, N1115);
not NOT1 (N2720, N2704);
buf BUF1 (N2721, N2719);
nor NOR4 (N2722, N2703, N684, N1635, N1247);
nand NAND4 (N2723, N2717, N1351, N1066, N653);
not NOT1 (N2724, N2711);
or OR2 (N2725, N2713, N2006);
not NOT1 (N2726, N2716);
not NOT1 (N2727, N2723);
nand NAND3 (N2728, N2724, N1435, N658);
nor NOR2 (N2729, N2725, N1010);
nand NAND2 (N2730, N2718, N90);
or OR3 (N2731, N2730, N1504, N683);
or OR4 (N2732, N2727, N964, N88, N2326);
nor NOR4 (N2733, N2731, N1479, N1931, N1253);
nand NAND4 (N2734, N2728, N2307, N1245, N2612);
or OR2 (N2735, N2729, N1170);
not NOT1 (N2736, N2735);
or OR3 (N2737, N2721, N1773, N1609);
or OR3 (N2738, N2734, N1136, N2477);
nor NOR4 (N2739, N2732, N250, N2439, N323);
not NOT1 (N2740, N2726);
nor NOR2 (N2741, N2737, N579);
and AND3 (N2742, N2706, N1955, N109);
not NOT1 (N2743, N2733);
nor NOR2 (N2744, N2715, N578);
xor XOR2 (N2745, N2738, N829);
xor XOR2 (N2746, N2742, N1369);
nand NAND3 (N2747, N2736, N2553, N232);
not NOT1 (N2748, N2747);
and AND2 (N2749, N2720, N1326);
not NOT1 (N2750, N2740);
and AND3 (N2751, N2743, N1776, N1702);
xor XOR2 (N2752, N2722, N1129);
buf BUF1 (N2753, N2751);
or OR2 (N2754, N2749, N7);
not NOT1 (N2755, N2741);
and AND2 (N2756, N2744, N391);
xor XOR2 (N2757, N2745, N144);
nor NOR2 (N2758, N2752, N1911);
nand NAND2 (N2759, N2754, N2291);
and AND2 (N2760, N2746, N2216);
or OR2 (N2761, N2759, N1065);
xor XOR2 (N2762, N2753, N1898);
not NOT1 (N2763, N2756);
or OR2 (N2764, N2750, N547);
xor XOR2 (N2765, N2764, N1719);
nor NOR4 (N2766, N2758, N519, N41, N2359);
buf BUF1 (N2767, N2755);
xor XOR2 (N2768, N2765, N1102);
not NOT1 (N2769, N2760);
nor NOR3 (N2770, N2768, N370, N1917);
xor XOR2 (N2771, N2767, N3);
nand NAND2 (N2772, N2757, N981);
or OR3 (N2773, N2739, N635, N941);
not NOT1 (N2774, N2748);
nor NOR4 (N2775, N2762, N256, N106, N2372);
or OR2 (N2776, N2774, N656);
buf BUF1 (N2777, N2771);
nor NOR2 (N2778, N2766, N294);
or OR2 (N2779, N2777, N1328);
nor NOR2 (N2780, N2775, N1565);
not NOT1 (N2781, N2769);
or OR2 (N2782, N2770, N1520);
and AND4 (N2783, N2761, N454, N2328, N1428);
nand NAND3 (N2784, N2778, N1586, N1638);
and AND3 (N2785, N2773, N1559, N1213);
nor NOR2 (N2786, N2779, N1365);
not NOT1 (N2787, N2784);
and AND3 (N2788, N2776, N1319, N2151);
nand NAND4 (N2789, N2782, N1990, N2606, N1380);
not NOT1 (N2790, N2788);
or OR2 (N2791, N2789, N698);
nor NOR4 (N2792, N2772, N2318, N2658, N2265);
or OR4 (N2793, N2763, N1222, N832, N645);
nor NOR2 (N2794, N2783, N663);
nand NAND3 (N2795, N2794, N2106, N386);
or OR4 (N2796, N2791, N1043, N77, N1950);
nor NOR2 (N2797, N2793, N1113);
nand NAND2 (N2798, N2795, N9);
or OR2 (N2799, N2790, N516);
nor NOR3 (N2800, N2799, N427, N828);
and AND4 (N2801, N2797, N2295, N162, N1445);
xor XOR2 (N2802, N2801, N752);
xor XOR2 (N2803, N2802, N319);
buf BUF1 (N2804, N2796);
and AND3 (N2805, N2785, N451, N762);
nand NAND4 (N2806, N2781, N1665, N623, N2743);
buf BUF1 (N2807, N2805);
and AND2 (N2808, N2798, N1776);
xor XOR2 (N2809, N2786, N2204);
or OR4 (N2810, N2804, N944, N1684, N1615);
xor XOR2 (N2811, N2809, N2346);
nand NAND3 (N2812, N2780, N2041, N130);
or OR3 (N2813, N2811, N1183, N1125);
and AND3 (N2814, N2787, N310, N1306);
and AND3 (N2815, N2803, N1257, N1570);
nor NOR2 (N2816, N2792, N483);
nor NOR4 (N2817, N2810, N2559, N2679, N1436);
nor NOR3 (N2818, N2817, N1053, N2381);
buf BUF1 (N2819, N2808);
buf BUF1 (N2820, N2807);
buf BUF1 (N2821, N2818);
or OR2 (N2822, N2816, N170);
and AND2 (N2823, N2815, N1486);
or OR4 (N2824, N2821, N1063, N2552, N2449);
nor NOR2 (N2825, N2823, N1347);
nor NOR3 (N2826, N2800, N2322, N2684);
nand NAND2 (N2827, N2824, N2480);
or OR3 (N2828, N2814, N1704, N2759);
buf BUF1 (N2829, N2825);
nor NOR3 (N2830, N2813, N2374, N645);
xor XOR2 (N2831, N2806, N1899);
or OR2 (N2832, N2812, N1296);
nand NAND4 (N2833, N2829, N1186, N983, N1505);
not NOT1 (N2834, N2833);
nor NOR4 (N2835, N2822, N2307, N88, N2120);
buf BUF1 (N2836, N2828);
buf BUF1 (N2837, N2834);
buf BUF1 (N2838, N2819);
buf BUF1 (N2839, N2831);
nor NOR3 (N2840, N2832, N816, N237);
nand NAND3 (N2841, N2835, N82, N1646);
buf BUF1 (N2842, N2827);
xor XOR2 (N2843, N2839, N2132);
not NOT1 (N2844, N2837);
nand NAND3 (N2845, N2842, N2808, N2153);
not NOT1 (N2846, N2845);
buf BUF1 (N2847, N2820);
buf BUF1 (N2848, N2844);
xor XOR2 (N2849, N2848, N859);
not NOT1 (N2850, N2841);
buf BUF1 (N2851, N2843);
nand NAND3 (N2852, N2826, N2414, N1291);
nor NOR4 (N2853, N2838, N779, N2625, N1294);
and AND3 (N2854, N2830, N2037, N1785);
not NOT1 (N2855, N2840);
and AND4 (N2856, N2855, N318, N2152, N856);
and AND2 (N2857, N2850, N1713);
nor NOR3 (N2858, N2847, N787, N1789);
buf BUF1 (N2859, N2836);
or OR2 (N2860, N2854, N2244);
buf BUF1 (N2861, N2856);
nor NOR3 (N2862, N2853, N2277, N1755);
and AND2 (N2863, N2849, N360);
and AND4 (N2864, N2861, N2807, N2631, N1997);
or OR3 (N2865, N2858, N2503, N502);
nor NOR4 (N2866, N2864, N1336, N2703, N1635);
buf BUF1 (N2867, N2863);
nor NOR2 (N2868, N2859, N313);
nand NAND4 (N2869, N2862, N2764, N246, N69);
xor XOR2 (N2870, N2869, N1763);
and AND2 (N2871, N2857, N537);
not NOT1 (N2872, N2867);
not NOT1 (N2873, N2870);
xor XOR2 (N2874, N2865, N2006);
xor XOR2 (N2875, N2871, N1738);
buf BUF1 (N2876, N2860);
and AND3 (N2877, N2873, N694, N2648);
buf BUF1 (N2878, N2876);
buf BUF1 (N2879, N2872);
or OR3 (N2880, N2846, N246, N1844);
buf BUF1 (N2881, N2880);
not NOT1 (N2882, N2877);
nor NOR3 (N2883, N2879, N655, N2546);
buf BUF1 (N2884, N2878);
xor XOR2 (N2885, N2851, N1471);
or OR4 (N2886, N2881, N403, N1278, N650);
or OR2 (N2887, N2868, N1022);
buf BUF1 (N2888, N2882);
nor NOR4 (N2889, N2883, N2771, N1285, N1548);
nor NOR2 (N2890, N2889, N1371);
xor XOR2 (N2891, N2888, N2845);
nand NAND3 (N2892, N2886, N2161, N583);
not NOT1 (N2893, N2874);
buf BUF1 (N2894, N2892);
or OR2 (N2895, N2875, N2198);
or OR3 (N2896, N2884, N2859, N1100);
buf BUF1 (N2897, N2866);
not NOT1 (N2898, N2885);
buf BUF1 (N2899, N2898);
nand NAND3 (N2900, N2891, N2604, N318);
or OR3 (N2901, N2887, N1235, N1451);
not NOT1 (N2902, N2897);
and AND2 (N2903, N2890, N365);
and AND3 (N2904, N2893, N1996, N66);
nand NAND4 (N2905, N2894, N864, N1655, N387);
not NOT1 (N2906, N2905);
buf BUF1 (N2907, N2903);
or OR3 (N2908, N2900, N2321, N2513);
or OR2 (N2909, N2906, N66);
nor NOR4 (N2910, N2852, N2411, N1844, N2510);
nor NOR2 (N2911, N2908, N1650);
nor NOR3 (N2912, N2899, N2238, N2365);
and AND4 (N2913, N2901, N1855, N1040, N571);
buf BUF1 (N2914, N2896);
not NOT1 (N2915, N2912);
or OR2 (N2916, N2911, N672);
not NOT1 (N2917, N2915);
nand NAND3 (N2918, N2909, N1934, N527);
nand NAND4 (N2919, N2904, N193, N718, N1537);
and AND3 (N2920, N2907, N422, N2389);
nor NOR2 (N2921, N2918, N2874);
not NOT1 (N2922, N2910);
not NOT1 (N2923, N2914);
nor NOR4 (N2924, N2920, N227, N405, N2712);
and AND4 (N2925, N2902, N2882, N302, N935);
nor NOR2 (N2926, N2919, N312);
not NOT1 (N2927, N2922);
xor XOR2 (N2928, N2923, N939);
xor XOR2 (N2929, N2921, N2252);
or OR3 (N2930, N2913, N85, N1019);
buf BUF1 (N2931, N2927);
not NOT1 (N2932, N2916);
xor XOR2 (N2933, N2926, N1625);
nor NOR4 (N2934, N2929, N1893, N67, N1319);
buf BUF1 (N2935, N2934);
and AND2 (N2936, N2924, N1276);
xor XOR2 (N2937, N2933, N2044);
xor XOR2 (N2938, N2935, N1649);
xor XOR2 (N2939, N2937, N1303);
not NOT1 (N2940, N2928);
nand NAND3 (N2941, N2925, N2746, N52);
not NOT1 (N2942, N2941);
xor XOR2 (N2943, N2930, N1094);
nor NOR4 (N2944, N2942, N1225, N2611, N1769);
or OR3 (N2945, N2932, N963, N2899);
xor XOR2 (N2946, N2940, N273);
xor XOR2 (N2947, N2945, N840);
and AND4 (N2948, N2943, N302, N1573, N2852);
buf BUF1 (N2949, N2948);
nor NOR2 (N2950, N2936, N124);
and AND2 (N2951, N2950, N1974);
buf BUF1 (N2952, N2947);
buf BUF1 (N2953, N2949);
buf BUF1 (N2954, N2953);
buf BUF1 (N2955, N2944);
nand NAND3 (N2956, N2939, N2040, N2436);
or OR3 (N2957, N2895, N2450, N1503);
and AND2 (N2958, N2917, N1330);
and AND3 (N2959, N2958, N2400, N1987);
not NOT1 (N2960, N2931);
not NOT1 (N2961, N2959);
or OR2 (N2962, N2955, N996);
xor XOR2 (N2963, N2952, N1138);
nand NAND4 (N2964, N2960, N394, N454, N1681);
nor NOR4 (N2965, N2954, N2297, N2927, N1217);
or OR2 (N2966, N2938, N2957);
not NOT1 (N2967, N2654);
xor XOR2 (N2968, N2951, N1790);
not NOT1 (N2969, N2963);
and AND4 (N2970, N2968, N1606, N1928, N128);
buf BUF1 (N2971, N2962);
xor XOR2 (N2972, N2956, N97);
nor NOR3 (N2973, N2970, N760, N668);
buf BUF1 (N2974, N2969);
nor NOR3 (N2975, N2965, N2336, N2109);
buf BUF1 (N2976, N2967);
or OR3 (N2977, N2974, N1658, N2385);
not NOT1 (N2978, N2976);
buf BUF1 (N2979, N2971);
or OR3 (N2980, N2973, N2587, N1515);
nand NAND3 (N2981, N2980, N1709, N1339);
xor XOR2 (N2982, N2977, N1542);
not NOT1 (N2983, N2966);
not NOT1 (N2984, N2979);
and AND2 (N2985, N2964, N2300);
nor NOR3 (N2986, N2984, N255, N485);
nor NOR3 (N2987, N2986, N1847, N2549);
or OR3 (N2988, N2983, N1938, N2153);
buf BUF1 (N2989, N2982);
nor NOR3 (N2990, N2989, N1216, N277);
not NOT1 (N2991, N2978);
xor XOR2 (N2992, N2991, N2167);
not NOT1 (N2993, N2981);
nand NAND4 (N2994, N2946, N2941, N1384, N501);
nor NOR4 (N2995, N2992, N2518, N2188, N2926);
not NOT1 (N2996, N2993);
or OR3 (N2997, N2996, N706, N1695);
xor XOR2 (N2998, N2975, N2188);
nor NOR4 (N2999, N2985, N1418, N2137, N1958);
not NOT1 (N3000, N2990);
nor NOR3 (N3001, N2998, N1391, N168);
xor XOR2 (N3002, N3000, N1923);
xor XOR2 (N3003, N2997, N2608);
nand NAND4 (N3004, N3003, N295, N2773, N911);
not NOT1 (N3005, N3002);
xor XOR2 (N3006, N2994, N2473);
not NOT1 (N3007, N3006);
and AND4 (N3008, N2988, N2671, N2981, N989);
not NOT1 (N3009, N3008);
nand NAND4 (N3010, N2987, N1980, N392, N1302);
and AND2 (N3011, N3007, N730);
xor XOR2 (N3012, N3001, N938);
and AND3 (N3013, N3012, N992, N1554);
or OR4 (N3014, N2961, N1697, N2392, N1430);
nand NAND2 (N3015, N2972, N2999);
nor NOR4 (N3016, N259, N1060, N1835, N55);
nand NAND3 (N3017, N3004, N2003, N629);
not NOT1 (N3018, N3015);
nand NAND4 (N3019, N3011, N1010, N1812, N360);
nand NAND2 (N3020, N3009, N3002);
nand NAND4 (N3021, N3019, N2824, N2787, N413);
nand NAND2 (N3022, N3021, N2998);
not NOT1 (N3023, N3005);
nor NOR2 (N3024, N3013, N425);
not NOT1 (N3025, N3010);
not NOT1 (N3026, N2995);
xor XOR2 (N3027, N3014, N2023);
or OR4 (N3028, N3024, N2257, N1435, N1349);
not NOT1 (N3029, N3027);
or OR2 (N3030, N3026, N490);
nor NOR2 (N3031, N3025, N1913);
nor NOR2 (N3032, N3020, N544);
nor NOR3 (N3033, N3022, N564, N913);
or OR2 (N3034, N3032, N1539);
or OR4 (N3035, N3029, N1090, N2396, N840);
not NOT1 (N3036, N3016);
buf BUF1 (N3037, N3033);
nand NAND4 (N3038, N3030, N2217, N2493, N2252);
buf BUF1 (N3039, N3036);
buf BUF1 (N3040, N3039);
or OR4 (N3041, N3017, N409, N1069, N2985);
nand NAND2 (N3042, N3040, N2725);
nor NOR4 (N3043, N3042, N1512, N220, N1359);
xor XOR2 (N3044, N3037, N1901);
nand NAND4 (N3045, N3031, N1397, N1083, N1119);
not NOT1 (N3046, N3023);
nand NAND3 (N3047, N3034, N2859, N1260);
nor NOR4 (N3048, N3028, N2324, N768, N2511);
nor NOR4 (N3049, N3043, N791, N490, N1497);
buf BUF1 (N3050, N3045);
and AND3 (N3051, N3038, N836, N1475);
nand NAND4 (N3052, N3041, N1768, N797, N2778);
xor XOR2 (N3053, N3044, N1068);
and AND3 (N3054, N3048, N1447, N1367);
or OR3 (N3055, N3053, N808, N1308);
xor XOR2 (N3056, N3047, N1864);
nand NAND4 (N3057, N3052, N784, N1207, N575);
not NOT1 (N3058, N3018);
and AND3 (N3059, N3054, N2840, N1209);
nand NAND4 (N3060, N3055, N2206, N2526, N3058);
buf BUF1 (N3061, N2905);
or OR4 (N3062, N3059, N2073, N1782, N385);
nand NAND2 (N3063, N3051, N2195);
not NOT1 (N3064, N3050);
and AND3 (N3065, N3056, N2083, N2586);
xor XOR2 (N3066, N3065, N1787);
not NOT1 (N3067, N3035);
and AND4 (N3068, N3060, N2215, N1223, N2580);
nand NAND3 (N3069, N3061, N1506, N1975);
and AND3 (N3070, N3057, N794, N2606);
buf BUF1 (N3071, N3067);
or OR4 (N3072, N3062, N1319, N641, N1233);
nor NOR4 (N3073, N3064, N383, N2933, N2381);
xor XOR2 (N3074, N3049, N924);
and AND3 (N3075, N3063, N2494, N230);
buf BUF1 (N3076, N3070);
or OR4 (N3077, N3046, N2, N2205, N1428);
nand NAND3 (N3078, N3068, N2086, N1019);
xor XOR2 (N3079, N3072, N217);
buf BUF1 (N3080, N3071);
nand NAND2 (N3081, N3076, N999);
xor XOR2 (N3082, N3079, N1126);
xor XOR2 (N3083, N3080, N1432);
xor XOR2 (N3084, N3066, N1919);
or OR2 (N3085, N3082, N1752);
nand NAND3 (N3086, N3078, N737, N2946);
nand NAND4 (N3087, N3085, N2437, N2098, N2169);
or OR3 (N3088, N3086, N84, N2341);
not NOT1 (N3089, N3088);
buf BUF1 (N3090, N3089);
or OR4 (N3091, N3075, N1260, N310, N629);
nand NAND2 (N3092, N3073, N363);
not NOT1 (N3093, N3074);
nand NAND2 (N3094, N3081, N1778);
xor XOR2 (N3095, N3090, N7);
and AND4 (N3096, N3093, N1786, N1350, N995);
xor XOR2 (N3097, N3087, N1488);
buf BUF1 (N3098, N3083);
not NOT1 (N3099, N3091);
or OR3 (N3100, N3092, N2990, N1045);
nand NAND3 (N3101, N3099, N1755, N267);
not NOT1 (N3102, N3069);
nor NOR3 (N3103, N3077, N3089, N1263);
nor NOR3 (N3104, N3095, N1004, N2876);
buf BUF1 (N3105, N3102);
or OR2 (N3106, N3104, N244);
xor XOR2 (N3107, N3105, N568);
and AND2 (N3108, N3103, N2725);
buf BUF1 (N3109, N3100);
not NOT1 (N3110, N3107);
nand NAND3 (N3111, N3084, N1775, N1978);
and AND4 (N3112, N3109, N525, N2182, N332);
and AND3 (N3113, N3110, N2729, N898);
not NOT1 (N3114, N3096);
or OR3 (N3115, N3113, N1340, N2660);
nor NOR4 (N3116, N3112, N2020, N463, N1756);
and AND4 (N3117, N3114, N2409, N2136, N2929);
buf BUF1 (N3118, N3098);
nor NOR4 (N3119, N3117, N1390, N425, N1694);
not NOT1 (N3120, N3101);
xor XOR2 (N3121, N3097, N2651);
nor NOR4 (N3122, N3121, N2864, N2825, N1792);
and AND4 (N3123, N3106, N2301, N2122, N2903);
or OR2 (N3124, N3108, N1871);
nand NAND2 (N3125, N3115, N288);
not NOT1 (N3126, N3116);
nor NOR3 (N3127, N3122, N2233, N2551);
nor NOR4 (N3128, N3127, N69, N519, N1873);
or OR4 (N3129, N3126, N1118, N1612, N1627);
not NOT1 (N3130, N3120);
and AND3 (N3131, N3094, N2352, N115);
nand NAND4 (N3132, N3118, N1199, N3108, N1397);
and AND2 (N3133, N3123, N2450);
not NOT1 (N3134, N3119);
or OR3 (N3135, N3125, N1520, N1472);
and AND4 (N3136, N3130, N1378, N2565, N370);
nand NAND4 (N3137, N3134, N2395, N2581, N150);
nor NOR2 (N3138, N3136, N412);
not NOT1 (N3139, N3131);
buf BUF1 (N3140, N3128);
not NOT1 (N3141, N3132);
nor NOR2 (N3142, N3137, N543);
and AND3 (N3143, N3124, N1598, N559);
or OR4 (N3144, N3129, N2861, N2114, N2160);
buf BUF1 (N3145, N3138);
not NOT1 (N3146, N3142);
not NOT1 (N3147, N3146);
and AND4 (N3148, N3143, N2841, N1882, N1546);
buf BUF1 (N3149, N3147);
or OR2 (N3150, N3133, N3112);
or OR4 (N3151, N3150, N97, N2043, N2705);
xor XOR2 (N3152, N3140, N1356);
nand NAND3 (N3153, N3149, N969, N2552);
not NOT1 (N3154, N3144);
nand NAND3 (N3155, N3145, N797, N1144);
or OR4 (N3156, N3111, N1714, N1618, N2482);
nor NOR4 (N3157, N3154, N938, N1611, N1654);
xor XOR2 (N3158, N3139, N2805);
buf BUF1 (N3159, N3148);
nand NAND3 (N3160, N3155, N756, N1955);
nor NOR3 (N3161, N3156, N2955, N465);
not NOT1 (N3162, N3135);
or OR3 (N3163, N3160, N711, N2875);
xor XOR2 (N3164, N3153, N3007);
or OR3 (N3165, N3163, N1067, N213);
nand NAND4 (N3166, N3151, N1232, N1952, N1723);
buf BUF1 (N3167, N3141);
xor XOR2 (N3168, N3162, N729);
xor XOR2 (N3169, N3158, N657);
buf BUF1 (N3170, N3165);
nand NAND2 (N3171, N3159, N1385);
not NOT1 (N3172, N3157);
or OR4 (N3173, N3170, N256, N156, N2146);
or OR2 (N3174, N3161, N571);
buf BUF1 (N3175, N3171);
and AND2 (N3176, N3166, N914);
nand NAND4 (N3177, N3169, N1162, N418, N2481);
not NOT1 (N3178, N3167);
and AND2 (N3179, N3174, N2382);
xor XOR2 (N3180, N3173, N2853);
or OR2 (N3181, N3175, N1790);
xor XOR2 (N3182, N3179, N2734);
or OR3 (N3183, N3178, N1663, N569);
buf BUF1 (N3184, N3168);
nor NOR2 (N3185, N3183, N2222);
buf BUF1 (N3186, N3164);
or OR3 (N3187, N3181, N1148, N1673);
nor NOR3 (N3188, N3152, N2871, N2074);
not NOT1 (N3189, N3184);
nor NOR2 (N3190, N3186, N2876);
nor NOR3 (N3191, N3177, N3046, N1249);
or OR3 (N3192, N3191, N1413, N222);
xor XOR2 (N3193, N3189, N325);
and AND2 (N3194, N3187, N1834);
xor XOR2 (N3195, N3193, N3066);
not NOT1 (N3196, N3195);
xor XOR2 (N3197, N3194, N1839);
nand NAND3 (N3198, N3182, N2559, N940);
not NOT1 (N3199, N3172);
buf BUF1 (N3200, N3176);
not NOT1 (N3201, N3200);
or OR4 (N3202, N3198, N2411, N2495, N1901);
or OR3 (N3203, N3202, N2964, N2026);
not NOT1 (N3204, N3199);
xor XOR2 (N3205, N3204, N280);
and AND3 (N3206, N3201, N2809, N2767);
not NOT1 (N3207, N3205);
nor NOR4 (N3208, N3185, N2282, N2996, N1507);
not NOT1 (N3209, N3197);
nand NAND3 (N3210, N3190, N1277, N1759);
buf BUF1 (N3211, N3208);
xor XOR2 (N3212, N3207, N111);
xor XOR2 (N3213, N3192, N2271);
xor XOR2 (N3214, N3209, N2261);
nor NOR4 (N3215, N3188, N3206, N2887, N2483);
not NOT1 (N3216, N3153);
nor NOR3 (N3217, N3211, N828, N909);
nor NOR2 (N3218, N3217, N2777);
not NOT1 (N3219, N3210);
xor XOR2 (N3220, N3219, N2083);
buf BUF1 (N3221, N3215);
nand NAND3 (N3222, N3212, N803, N2429);
nand NAND2 (N3223, N3222, N389);
nor NOR3 (N3224, N3213, N1077, N2007);
nand NAND2 (N3225, N3203, N581);
nand NAND4 (N3226, N3225, N2863, N1902, N625);
and AND3 (N3227, N3224, N2354, N1246);
nand NAND4 (N3228, N3180, N2205, N1372, N932);
not NOT1 (N3229, N3226);
not NOT1 (N3230, N3229);
nand NAND2 (N3231, N3223, N754);
xor XOR2 (N3232, N3220, N1374);
xor XOR2 (N3233, N3218, N2499);
nor NOR3 (N3234, N3228, N1755, N455);
xor XOR2 (N3235, N3234, N716);
nor NOR2 (N3236, N3231, N1135);
nand NAND2 (N3237, N3216, N2482);
or OR4 (N3238, N3230, N551, N2966, N1461);
nor NOR4 (N3239, N3232, N497, N2585, N374);
not NOT1 (N3240, N3221);
xor XOR2 (N3241, N3227, N814);
nand NAND3 (N3242, N3240, N2939, N749);
nand NAND3 (N3243, N3236, N1597, N1154);
xor XOR2 (N3244, N3196, N231);
or OR2 (N3245, N3241, N1764);
xor XOR2 (N3246, N3239, N308);
buf BUF1 (N3247, N3237);
and AND4 (N3248, N3235, N1385, N1274, N2143);
nand NAND2 (N3249, N3242, N1517);
nand NAND3 (N3250, N3244, N735, N90);
nand NAND4 (N3251, N3245, N1098, N1905, N2011);
nand NAND2 (N3252, N3214, N601);
or OR4 (N3253, N3243, N1799, N2390, N2420);
and AND4 (N3254, N3252, N1884, N1235, N2919);
nor NOR3 (N3255, N3238, N263, N1207);
or OR4 (N3256, N3251, N1999, N722, N695);
nand NAND3 (N3257, N3248, N1119, N1158);
nand NAND3 (N3258, N3254, N480, N209);
or OR4 (N3259, N3253, N880, N2458, N2393);
xor XOR2 (N3260, N3256, N1875);
or OR2 (N3261, N3246, N1928);
buf BUF1 (N3262, N3258);
buf BUF1 (N3263, N3247);
not NOT1 (N3264, N3255);
not NOT1 (N3265, N3250);
not NOT1 (N3266, N3233);
buf BUF1 (N3267, N3257);
and AND3 (N3268, N3262, N2512, N2819);
or OR4 (N3269, N3261, N2608, N2843, N2089);
and AND2 (N3270, N3268, N1502);
nor NOR4 (N3271, N3270, N816, N2487, N1832);
and AND4 (N3272, N3271, N1823, N466, N2245);
xor XOR2 (N3273, N3264, N2576);
buf BUF1 (N3274, N3273);
and AND2 (N3275, N3269, N1304);
not NOT1 (N3276, N3274);
nor NOR3 (N3277, N3259, N251, N1288);
and AND2 (N3278, N3266, N796);
nand NAND3 (N3279, N3267, N983, N681);
and AND3 (N3280, N3278, N1447, N1667);
not NOT1 (N3281, N3260);
and AND3 (N3282, N3279, N1638, N1057);
or OR2 (N3283, N3272, N2226);
not NOT1 (N3284, N3249);
not NOT1 (N3285, N3265);
and AND4 (N3286, N3263, N2463, N592, N1411);
buf BUF1 (N3287, N3284);
nor NOR3 (N3288, N3282, N2944, N768);
xor XOR2 (N3289, N3286, N889);
nor NOR2 (N3290, N3277, N160);
not NOT1 (N3291, N3281);
nand NAND2 (N3292, N3291, N2414);
buf BUF1 (N3293, N3283);
nor NOR3 (N3294, N3276, N558, N1068);
nand NAND3 (N3295, N3294, N1836, N1943);
nor NOR3 (N3296, N3289, N137, N957);
or OR4 (N3297, N3280, N1341, N2664, N1569);
nand NAND3 (N3298, N3290, N1970, N567);
buf BUF1 (N3299, N3285);
nand NAND3 (N3300, N3288, N1388, N473);
nor NOR4 (N3301, N3292, N2303, N567, N465);
xor XOR2 (N3302, N3300, N192);
not NOT1 (N3303, N3298);
or OR4 (N3304, N3299, N678, N1190, N1844);
buf BUF1 (N3305, N3304);
nand NAND4 (N3306, N3296, N1775, N2777, N2422);
not NOT1 (N3307, N3301);
nor NOR3 (N3308, N3302, N1461, N1350);
or OR4 (N3309, N3295, N2375, N1300, N681);
and AND4 (N3310, N3308, N1341, N1326, N2928);
nand NAND2 (N3311, N3309, N2091);
not NOT1 (N3312, N3287);
buf BUF1 (N3313, N3303);
and AND2 (N3314, N3312, N2211);
buf BUF1 (N3315, N3293);
xor XOR2 (N3316, N3307, N2784);
and AND3 (N3317, N3306, N551, N980);
nor NOR4 (N3318, N3297, N2166, N3288, N448);
xor XOR2 (N3319, N3305, N2490);
nor NOR3 (N3320, N3310, N2328, N288);
nand NAND3 (N3321, N3275, N626, N3288);
xor XOR2 (N3322, N3317, N1689);
nand NAND2 (N3323, N3319, N3010);
and AND3 (N3324, N3320, N1339, N1456);
buf BUF1 (N3325, N3322);
and AND4 (N3326, N3318, N3232, N2123, N1311);
xor XOR2 (N3327, N3316, N2727);
and AND3 (N3328, N3326, N2351, N1709);
xor XOR2 (N3329, N3314, N467);
or OR2 (N3330, N3323, N2925);
nand NAND3 (N3331, N3313, N75, N1991);
buf BUF1 (N3332, N3324);
nor NOR3 (N3333, N3328, N504, N1751);
or OR2 (N3334, N3311, N3274);
and AND2 (N3335, N3315, N2069);
and AND2 (N3336, N3325, N1003);
or OR4 (N3337, N3336, N1398, N823, N3012);
nand NAND4 (N3338, N3327, N2897, N3119, N1263);
or OR2 (N3339, N3332, N1428);
or OR4 (N3340, N3338, N2459, N3108, N1384);
or OR2 (N3341, N3337, N3147);
nand NAND4 (N3342, N3339, N1879, N1337, N1674);
or OR4 (N3343, N3341, N315, N3255, N2986);
or OR2 (N3344, N3321, N2589);
nand NAND4 (N3345, N3333, N907, N2571, N717);
nor NOR4 (N3346, N3331, N2431, N1764, N2370);
or OR4 (N3347, N3344, N838, N2686, N2738);
nor NOR2 (N3348, N3345, N1076);
and AND3 (N3349, N3347, N602, N2062);
and AND3 (N3350, N3346, N1380, N2034);
xor XOR2 (N3351, N3340, N1009);
xor XOR2 (N3352, N3330, N471);
nand NAND2 (N3353, N3350, N2980);
nand NAND4 (N3354, N3335, N2310, N997, N2937);
buf BUF1 (N3355, N3353);
nor NOR2 (N3356, N3354, N2085);
nor NOR2 (N3357, N3348, N1727);
not NOT1 (N3358, N3343);
nand NAND2 (N3359, N3342, N817);
xor XOR2 (N3360, N3355, N757);
or OR4 (N3361, N3352, N208, N1112, N2080);
buf BUF1 (N3362, N3360);
xor XOR2 (N3363, N3357, N975);
xor XOR2 (N3364, N3363, N1859);
nand NAND3 (N3365, N3351, N2516, N2714);
buf BUF1 (N3366, N3365);
xor XOR2 (N3367, N3329, N1296);
or OR3 (N3368, N3361, N669, N2);
buf BUF1 (N3369, N3358);
nand NAND2 (N3370, N3367, N822);
nand NAND3 (N3371, N3366, N149, N327);
buf BUF1 (N3372, N3359);
xor XOR2 (N3373, N3370, N3309);
nor NOR4 (N3374, N3362, N1390, N2311, N841);
not NOT1 (N3375, N3373);
buf BUF1 (N3376, N3375);
or OR4 (N3377, N3371, N86, N1741, N71);
nand NAND4 (N3378, N3372, N1084, N2964, N767);
not NOT1 (N3379, N3374);
xor XOR2 (N3380, N3334, N2862);
not NOT1 (N3381, N3356);
and AND3 (N3382, N3369, N1882, N1742);
xor XOR2 (N3383, N3381, N2674);
xor XOR2 (N3384, N3383, N2160);
or OR2 (N3385, N3349, N519);
buf BUF1 (N3386, N3368);
or OR2 (N3387, N3376, N3031);
or OR2 (N3388, N3380, N210);
nor NOR4 (N3389, N3384, N1952, N2912, N877);
buf BUF1 (N3390, N3382);
or OR2 (N3391, N3390, N608);
nor NOR3 (N3392, N3378, N1152, N699);
and AND4 (N3393, N3387, N1597, N1911, N3252);
xor XOR2 (N3394, N3389, N1005);
or OR4 (N3395, N3379, N3049, N37, N259);
and AND2 (N3396, N3393, N1788);
buf BUF1 (N3397, N3377);
not NOT1 (N3398, N3397);
not NOT1 (N3399, N3395);
not NOT1 (N3400, N3396);
not NOT1 (N3401, N3399);
nor NOR2 (N3402, N3385, N3142);
buf BUF1 (N3403, N3398);
or OR2 (N3404, N3400, N1548);
buf BUF1 (N3405, N3388);
not NOT1 (N3406, N3364);
not NOT1 (N3407, N3406);
or OR4 (N3408, N3405, N3278, N2303, N1407);
or OR4 (N3409, N3403, N1706, N849, N2823);
buf BUF1 (N3410, N3407);
and AND3 (N3411, N3401, N1312, N2086);
nor NOR2 (N3412, N3409, N898);
not NOT1 (N3413, N3408);
nand NAND3 (N3414, N3413, N596, N1855);
nor NOR4 (N3415, N3386, N3100, N304, N1279);
and AND3 (N3416, N3394, N3264, N996);
xor XOR2 (N3417, N3402, N3186);
buf BUF1 (N3418, N3417);
nand NAND2 (N3419, N3391, N907);
or OR3 (N3420, N3414, N1823, N1517);
buf BUF1 (N3421, N3410);
not NOT1 (N3422, N3415);
nand NAND4 (N3423, N3392, N1259, N3124, N651);
nor NOR2 (N3424, N3412, N506);
xor XOR2 (N3425, N3424, N3241);
nor NOR2 (N3426, N3404, N2752);
not NOT1 (N3427, N3416);
buf BUF1 (N3428, N3422);
nor NOR2 (N3429, N3426, N2591);
xor XOR2 (N3430, N3421, N2390);
or OR3 (N3431, N3423, N281, N550);
nand NAND2 (N3432, N3425, N1315);
buf BUF1 (N3433, N3418);
xor XOR2 (N3434, N3430, N1861);
not NOT1 (N3435, N3427);
and AND2 (N3436, N3431, N1964);
nor NOR3 (N3437, N3428, N647, N2673);
xor XOR2 (N3438, N3433, N1669);
nand NAND2 (N3439, N3419, N296);
and AND3 (N3440, N3439, N2151, N2003);
xor XOR2 (N3441, N3432, N263);
nor NOR3 (N3442, N3411, N230, N878);
buf BUF1 (N3443, N3441);
not NOT1 (N3444, N3440);
and AND4 (N3445, N3437, N943, N562, N321);
nor NOR4 (N3446, N3444, N1183, N1096, N2973);
xor XOR2 (N3447, N3445, N1329);
nor NOR4 (N3448, N3420, N2266, N3100, N2955);
xor XOR2 (N3449, N3448, N1154);
buf BUF1 (N3450, N3436);
nand NAND4 (N3451, N3434, N1478, N758, N501);
nand NAND2 (N3452, N3438, N701);
and AND4 (N3453, N3449, N3100, N1423, N2614);
and AND3 (N3454, N3435, N3450, N2032);
buf BUF1 (N3455, N2966);
not NOT1 (N3456, N3443);
and AND3 (N3457, N3454, N1334, N3109);
xor XOR2 (N3458, N3451, N1107);
or OR4 (N3459, N3453, N2085, N465, N453);
nand NAND3 (N3460, N3447, N2224, N2589);
not NOT1 (N3461, N3442);
buf BUF1 (N3462, N3456);
not NOT1 (N3463, N3458);
not NOT1 (N3464, N3461);
or OR4 (N3465, N3429, N928, N1759, N2066);
nor NOR2 (N3466, N3459, N199);
xor XOR2 (N3467, N3465, N2091);
nor NOR3 (N3468, N3466, N245, N3405);
xor XOR2 (N3469, N3455, N3228);
or OR3 (N3470, N3469, N1943, N1796);
and AND3 (N3471, N3468, N450, N37);
not NOT1 (N3472, N3463);
and AND4 (N3473, N3464, N526, N2943, N1634);
not NOT1 (N3474, N3472);
nand NAND2 (N3475, N3452, N494);
or OR4 (N3476, N3467, N1042, N1470, N1311);
nor NOR3 (N3477, N3474, N1191, N477);
nor NOR4 (N3478, N3446, N2373, N2809, N1503);
nand NAND3 (N3479, N3462, N1775, N33);
nor NOR3 (N3480, N3471, N400, N520);
not NOT1 (N3481, N3476);
not NOT1 (N3482, N3480);
not NOT1 (N3483, N3482);
xor XOR2 (N3484, N3477, N2913);
xor XOR2 (N3485, N3481, N975);
not NOT1 (N3486, N3484);
nor NOR2 (N3487, N3475, N3237);
not NOT1 (N3488, N3486);
and AND3 (N3489, N3473, N290, N2837);
or OR4 (N3490, N3485, N1124, N774, N268);
or OR3 (N3491, N3460, N2954, N596);
and AND2 (N3492, N3490, N3369);
not NOT1 (N3493, N3488);
and AND3 (N3494, N3487, N3266, N3276);
and AND2 (N3495, N3491, N1273);
nand NAND2 (N3496, N3470, N926);
not NOT1 (N3497, N3495);
or OR4 (N3498, N3497, N2945, N428, N806);
and AND4 (N3499, N3483, N2353, N3160, N2642);
buf BUF1 (N3500, N3492);
nand NAND2 (N3501, N3500, N898);
not NOT1 (N3502, N3494);
and AND4 (N3503, N3478, N2693, N951, N97);
buf BUF1 (N3504, N3489);
buf BUF1 (N3505, N3504);
xor XOR2 (N3506, N3457, N2279);
nor NOR4 (N3507, N3498, N1205, N1100, N1999);
xor XOR2 (N3508, N3501, N2952);
nor NOR2 (N3509, N3507, N2193);
nand NAND4 (N3510, N3496, N3425, N2225, N1337);
nor NOR2 (N3511, N3506, N713);
or OR3 (N3512, N3499, N3065, N540);
nand NAND2 (N3513, N3508, N55);
or OR4 (N3514, N3493, N1948, N2642, N1747);
or OR2 (N3515, N3513, N2484);
and AND2 (N3516, N3511, N2434);
or OR3 (N3517, N3510, N583, N2908);
and AND4 (N3518, N3503, N813, N546, N260);
buf BUF1 (N3519, N3505);
nand NAND2 (N3520, N3516, N3064);
not NOT1 (N3521, N3517);
nand NAND4 (N3522, N3521, N1902, N3450, N1799);
xor XOR2 (N3523, N3515, N1527);
xor XOR2 (N3524, N3519, N1107);
buf BUF1 (N3525, N3479);
nand NAND2 (N3526, N3514, N3223);
and AND4 (N3527, N3518, N1926, N3076, N1144);
xor XOR2 (N3528, N3523, N3187);
or OR3 (N3529, N3520, N1908, N1147);
or OR3 (N3530, N3528, N3465, N1023);
nor NOR2 (N3531, N3530, N1323);
xor XOR2 (N3532, N3502, N2288);
or OR2 (N3533, N3532, N709);
buf BUF1 (N3534, N3509);
nand NAND3 (N3535, N3533, N3352, N1093);
and AND2 (N3536, N3529, N1993);
and AND2 (N3537, N3536, N562);
buf BUF1 (N3538, N3524);
xor XOR2 (N3539, N3538, N2150);
nor NOR2 (N3540, N3535, N1168);
not NOT1 (N3541, N3537);
xor XOR2 (N3542, N3541, N1724);
not NOT1 (N3543, N3526);
buf BUF1 (N3544, N3534);
and AND3 (N3545, N3522, N1851, N1622);
and AND4 (N3546, N3543, N628, N1553, N113);
not NOT1 (N3547, N3525);
nand NAND4 (N3548, N3531, N404, N735, N1236);
xor XOR2 (N3549, N3542, N95);
buf BUF1 (N3550, N3512);
and AND4 (N3551, N3544, N2496, N930, N3085);
not NOT1 (N3552, N3545);
buf BUF1 (N3553, N3548);
and AND2 (N3554, N3551, N3098);
or OR3 (N3555, N3553, N342, N2302);
and AND3 (N3556, N3550, N626, N3418);
and AND3 (N3557, N3540, N1471, N541);
or OR3 (N3558, N3554, N3114, N442);
xor XOR2 (N3559, N3558, N420);
buf BUF1 (N3560, N3552);
nand NAND2 (N3561, N3560, N26);
nor NOR2 (N3562, N3527, N2829);
or OR2 (N3563, N3557, N3043);
and AND4 (N3564, N3539, N2746, N1962, N1729);
nor NOR3 (N3565, N3561, N908, N3483);
not NOT1 (N3566, N3564);
nor NOR4 (N3567, N3562, N1696, N1418, N2957);
nor NOR3 (N3568, N3546, N1272, N390);
not NOT1 (N3569, N3556);
or OR4 (N3570, N3568, N997, N1664, N2318);
xor XOR2 (N3571, N3547, N1131);
not NOT1 (N3572, N3549);
and AND2 (N3573, N3555, N617);
nor NOR4 (N3574, N3573, N3372, N2034, N793);
nor NOR2 (N3575, N3565, N2055);
not NOT1 (N3576, N3569);
buf BUF1 (N3577, N3566);
and AND3 (N3578, N3574, N640, N552);
xor XOR2 (N3579, N3572, N2661);
nor NOR4 (N3580, N3579, N409, N1113, N913);
nand NAND2 (N3581, N3576, N2453);
buf BUF1 (N3582, N3580);
buf BUF1 (N3583, N3582);
buf BUF1 (N3584, N3563);
nor NOR3 (N3585, N3575, N1343, N2335);
xor XOR2 (N3586, N3583, N2093);
buf BUF1 (N3587, N3578);
and AND4 (N3588, N3585, N2781, N198, N219);
xor XOR2 (N3589, N3588, N3151);
nand NAND2 (N3590, N3577, N3067);
nand NAND3 (N3591, N3584, N697, N3021);
or OR4 (N3592, N3571, N2170, N3534, N1156);
or OR2 (N3593, N3586, N2426);
and AND3 (N3594, N3567, N3334, N1145);
and AND2 (N3595, N3589, N3464);
and AND3 (N3596, N3559, N2818, N432);
nand NAND2 (N3597, N3590, N2144);
nand NAND3 (N3598, N3592, N774, N2536);
nand NAND2 (N3599, N3598, N1707);
xor XOR2 (N3600, N3587, N194);
and AND2 (N3601, N3595, N2813);
or OR3 (N3602, N3591, N3187, N605);
or OR3 (N3603, N3570, N253, N1864);
nor NOR2 (N3604, N3597, N2251);
not NOT1 (N3605, N3602);
and AND2 (N3606, N3604, N2066);
nand NAND4 (N3607, N3594, N2173, N562, N3522);
nor NOR3 (N3608, N3606, N1523, N2503);
and AND3 (N3609, N3593, N365, N184);
buf BUF1 (N3610, N3609);
buf BUF1 (N3611, N3610);
xor XOR2 (N3612, N3596, N3049);
nor NOR3 (N3613, N3601, N223, N336);
nand NAND2 (N3614, N3607, N572);
nor NOR4 (N3615, N3581, N1193, N11, N3586);
not NOT1 (N3616, N3614);
buf BUF1 (N3617, N3613);
not NOT1 (N3618, N3600);
xor XOR2 (N3619, N3599, N1808);
or OR3 (N3620, N3605, N2707, N1041);
not NOT1 (N3621, N3619);
buf BUF1 (N3622, N3611);
not NOT1 (N3623, N3620);
xor XOR2 (N3624, N3612, N3149);
xor XOR2 (N3625, N3618, N116);
buf BUF1 (N3626, N3616);
xor XOR2 (N3627, N3622, N2430);
and AND2 (N3628, N3623, N293);
or OR3 (N3629, N3621, N2485, N1259);
buf BUF1 (N3630, N3626);
nand NAND2 (N3631, N3617, N2278);
and AND2 (N3632, N3615, N3382);
nor NOR3 (N3633, N3627, N3249, N673);
and AND4 (N3634, N3608, N1457, N1955, N689);
nand NAND4 (N3635, N3631, N1560, N369, N1741);
nand NAND2 (N3636, N3632, N116);
or OR4 (N3637, N3630, N589, N1677, N2608);
not NOT1 (N3638, N3635);
buf BUF1 (N3639, N3634);
xor XOR2 (N3640, N3637, N783);
or OR4 (N3641, N3636, N917, N101, N192);
or OR2 (N3642, N3641, N998);
not NOT1 (N3643, N3628);
or OR3 (N3644, N3633, N2296, N203);
nor NOR3 (N3645, N3639, N2670, N3295);
not NOT1 (N3646, N3645);
not NOT1 (N3647, N3646);
buf BUF1 (N3648, N3629);
or OR3 (N3649, N3603, N3072, N2152);
buf BUF1 (N3650, N3638);
nand NAND2 (N3651, N3643, N3573);
buf BUF1 (N3652, N3650);
nand NAND4 (N3653, N3651, N268, N781, N1379);
nand NAND4 (N3654, N3648, N198, N258, N1536);
or OR4 (N3655, N3654, N2840, N1460, N406);
not NOT1 (N3656, N3655);
xor XOR2 (N3657, N3624, N1236);
xor XOR2 (N3658, N3656, N3377);
buf BUF1 (N3659, N3647);
or OR2 (N3660, N3659, N1742);
and AND3 (N3661, N3640, N2244, N2594);
nand NAND3 (N3662, N3649, N512, N1317);
or OR4 (N3663, N3642, N238, N443, N35);
buf BUF1 (N3664, N3660);
xor XOR2 (N3665, N3661, N1357);
nand NAND4 (N3666, N3662, N1882, N3594, N3036);
or OR2 (N3667, N3653, N1140);
buf BUF1 (N3668, N3666);
or OR3 (N3669, N3664, N1994, N889);
nor NOR2 (N3670, N3663, N419);
nand NAND3 (N3671, N3670, N746, N3403);
or OR4 (N3672, N3658, N255, N1803, N2542);
nand NAND3 (N3673, N3668, N597, N1072);
buf BUF1 (N3674, N3667);
buf BUF1 (N3675, N3665);
buf BUF1 (N3676, N3644);
buf BUF1 (N3677, N3657);
xor XOR2 (N3678, N3676, N2387);
or OR3 (N3679, N3652, N328, N199);
nor NOR3 (N3680, N3674, N3202, N1933);
nand NAND4 (N3681, N3673, N94, N2603, N2530);
not NOT1 (N3682, N3669);
and AND2 (N3683, N3682, N1800);
and AND4 (N3684, N3679, N3057, N2567, N3615);
or OR4 (N3685, N3625, N540, N3608, N2742);
nor NOR4 (N3686, N3685, N15, N1146, N2478);
not NOT1 (N3687, N3683);
or OR3 (N3688, N3675, N1895, N942);
and AND2 (N3689, N3671, N3387);
and AND2 (N3690, N3678, N970);
not NOT1 (N3691, N3686);
not NOT1 (N3692, N3689);
and AND3 (N3693, N3672, N948, N716);
or OR2 (N3694, N3680, N2747);
nor NOR4 (N3695, N3690, N957, N2836, N2248);
not NOT1 (N3696, N3691);
and AND4 (N3697, N3694, N294, N3029, N1895);
nand NAND2 (N3698, N3684, N2746);
xor XOR2 (N3699, N3677, N2797);
and AND4 (N3700, N3693, N1917, N67, N2881);
and AND2 (N3701, N3695, N3262);
or OR4 (N3702, N3700, N78, N1057, N3362);
xor XOR2 (N3703, N3698, N927);
nand NAND2 (N3704, N3697, N1201);
nand NAND2 (N3705, N3704, N2568);
nand NAND4 (N3706, N3702, N2043, N1857, N111);
nand NAND4 (N3707, N3705, N2951, N666, N3200);
buf BUF1 (N3708, N3681);
xor XOR2 (N3709, N3706, N159);
not NOT1 (N3710, N3701);
xor XOR2 (N3711, N3709, N2522);
not NOT1 (N3712, N3711);
not NOT1 (N3713, N3710);
xor XOR2 (N3714, N3712, N335);
or OR3 (N3715, N3688, N1412, N818);
nand NAND3 (N3716, N3713, N2395, N767);
buf BUF1 (N3717, N3714);
buf BUF1 (N3718, N3692);
nand NAND4 (N3719, N3717, N443, N1377, N1209);
xor XOR2 (N3720, N3687, N2554);
nor NOR3 (N3721, N3716, N651, N2336);
buf BUF1 (N3722, N3708);
nand NAND3 (N3723, N3719, N633, N2834);
and AND4 (N3724, N3707, N1178, N3077, N1593);
nand NAND2 (N3725, N3723, N3387);
not NOT1 (N3726, N3699);
and AND4 (N3727, N3721, N3536, N2388, N1480);
nand NAND3 (N3728, N3726, N1292, N152);
and AND3 (N3729, N3696, N3405, N2885);
not NOT1 (N3730, N3703);
and AND4 (N3731, N3727, N3106, N53, N134);
and AND3 (N3732, N3731, N705, N2889);
nor NOR3 (N3733, N3729, N3238, N1673);
xor XOR2 (N3734, N3722, N2405);
nand NAND3 (N3735, N3724, N3603, N3174);
nor NOR3 (N3736, N3733, N1372, N2168);
xor XOR2 (N3737, N3734, N2352);
nor NOR2 (N3738, N3715, N380);
and AND3 (N3739, N3718, N2790, N569);
nor NOR4 (N3740, N3738, N1068, N3022, N152);
or OR3 (N3741, N3739, N2630, N3581);
not NOT1 (N3742, N3730);
nor NOR3 (N3743, N3736, N1608, N1324);
nand NAND3 (N3744, N3742, N3155, N685);
not NOT1 (N3745, N3740);
and AND2 (N3746, N3737, N255);
not NOT1 (N3747, N3728);
nand NAND4 (N3748, N3732, N56, N2698, N2271);
or OR2 (N3749, N3720, N34);
nand NAND2 (N3750, N3748, N2902);
nand NAND3 (N3751, N3747, N1377, N1885);
not NOT1 (N3752, N3750);
or OR4 (N3753, N3743, N1241, N2144, N3032);
nand NAND4 (N3754, N3752, N369, N2152, N2118);
nand NAND4 (N3755, N3753, N1959, N572, N2647);
nand NAND4 (N3756, N3755, N203, N205, N3366);
or OR3 (N3757, N3744, N809, N648);
nor NOR2 (N3758, N3749, N1855);
and AND2 (N3759, N3746, N3669);
xor XOR2 (N3760, N3725, N805);
not NOT1 (N3761, N3760);
nand NAND2 (N3762, N3761, N1008);
buf BUF1 (N3763, N3762);
buf BUF1 (N3764, N3735);
and AND2 (N3765, N3763, N2026);
and AND3 (N3766, N3758, N730, N3759);
nand NAND3 (N3767, N1219, N3612, N2736);
or OR4 (N3768, N3765, N230, N1464, N3185);
or OR3 (N3769, N3756, N1445, N2888);
nand NAND3 (N3770, N3764, N1908, N3184);
nor NOR2 (N3771, N3754, N2405);
nand NAND2 (N3772, N3766, N3225);
nor NOR2 (N3773, N3770, N2836);
nand NAND3 (N3774, N3769, N1725, N3218);
buf BUF1 (N3775, N3741);
xor XOR2 (N3776, N3773, N2519);
nand NAND2 (N3777, N3768, N1022);
nand NAND2 (N3778, N3767, N3576);
or OR4 (N3779, N3745, N406, N2744, N3017);
not NOT1 (N3780, N3757);
or OR4 (N3781, N3776, N3158, N2233, N2835);
or OR3 (N3782, N3751, N117, N2141);
not NOT1 (N3783, N3774);
and AND2 (N3784, N3777, N1676);
and AND2 (N3785, N3771, N1054);
xor XOR2 (N3786, N3775, N1098);
not NOT1 (N3787, N3786);
nor NOR4 (N3788, N3781, N2526, N3248, N1082);
nand NAND3 (N3789, N3778, N3232, N371);
or OR3 (N3790, N3785, N1408, N2644);
or OR3 (N3791, N3787, N2424, N112);
and AND4 (N3792, N3788, N2014, N2108, N631);
buf BUF1 (N3793, N3791);
not NOT1 (N3794, N3784);
or OR3 (N3795, N3790, N2208, N3011);
xor XOR2 (N3796, N3772, N2427);
and AND2 (N3797, N3792, N1423);
xor XOR2 (N3798, N3795, N2614);
and AND3 (N3799, N3779, N2571, N2582);
or OR3 (N3800, N3782, N2163, N858);
nand NAND3 (N3801, N3798, N3354, N930);
nor NOR2 (N3802, N3801, N321);
and AND3 (N3803, N3796, N2399, N3058);
not NOT1 (N3804, N3794);
xor XOR2 (N3805, N3783, N3163);
and AND2 (N3806, N3805, N1896);
and AND3 (N3807, N3806, N1341, N1131);
and AND2 (N3808, N3803, N3704);
and AND3 (N3809, N3799, N1197, N1501);
and AND2 (N3810, N3797, N2936);
and AND2 (N3811, N3789, N3166);
buf BUF1 (N3812, N3802);
and AND4 (N3813, N3793, N3261, N2923, N2243);
xor XOR2 (N3814, N3810, N1324);
buf BUF1 (N3815, N3811);
or OR2 (N3816, N3808, N924);
not NOT1 (N3817, N3809);
not NOT1 (N3818, N3804);
not NOT1 (N3819, N3780);
nor NOR2 (N3820, N3812, N2835);
and AND3 (N3821, N3820, N2037, N3460);
and AND3 (N3822, N3818, N408, N521);
buf BUF1 (N3823, N3814);
xor XOR2 (N3824, N3822, N135);
nand NAND3 (N3825, N3824, N1685, N2033);
nand NAND2 (N3826, N3800, N3204);
xor XOR2 (N3827, N3817, N3219);
nor NOR2 (N3828, N3815, N1740);
not NOT1 (N3829, N3807);
nand NAND3 (N3830, N3816, N1302, N2201);
and AND2 (N3831, N3813, N913);
and AND2 (N3832, N3828, N2658);
and AND2 (N3833, N3831, N1640);
or OR4 (N3834, N3833, N765, N2186, N3166);
buf BUF1 (N3835, N3826);
xor XOR2 (N3836, N3830, N1639);
and AND4 (N3837, N3829, N1036, N2509, N438);
nor NOR3 (N3838, N3835, N422, N1731);
buf BUF1 (N3839, N3819);
and AND2 (N3840, N3834, N516);
not NOT1 (N3841, N3837);
xor XOR2 (N3842, N3823, N2729);
not NOT1 (N3843, N3832);
not NOT1 (N3844, N3839);
buf BUF1 (N3845, N3836);
nand NAND2 (N3846, N3838, N2141);
not NOT1 (N3847, N3845);
nand NAND2 (N3848, N3825, N751);
xor XOR2 (N3849, N3847, N2363);
buf BUF1 (N3850, N3840);
or OR2 (N3851, N3844, N1584);
nand NAND4 (N3852, N3848, N3109, N412, N2149);
not NOT1 (N3853, N3852);
xor XOR2 (N3854, N3849, N803);
nand NAND3 (N3855, N3827, N1712, N1727);
nor NOR3 (N3856, N3853, N99, N2364);
or OR2 (N3857, N3851, N118);
nand NAND3 (N3858, N3842, N772, N3801);
or OR3 (N3859, N3858, N3276, N231);
buf BUF1 (N3860, N3855);
buf BUF1 (N3861, N3841);
nor NOR2 (N3862, N3850, N2699);
not NOT1 (N3863, N3857);
not NOT1 (N3864, N3821);
nand NAND4 (N3865, N3859, N2753, N1193, N2675);
nand NAND3 (N3866, N3864, N193, N1746);
buf BUF1 (N3867, N3856);
nor NOR2 (N3868, N3865, N274);
and AND4 (N3869, N3846, N2131, N1756, N998);
nor NOR2 (N3870, N3868, N1742);
xor XOR2 (N3871, N3843, N793);
and AND4 (N3872, N3863, N2429, N2726, N674);
not NOT1 (N3873, N3862);
buf BUF1 (N3874, N3867);
xor XOR2 (N3875, N3872, N3643);
buf BUF1 (N3876, N3854);
or OR2 (N3877, N3861, N2736);
nand NAND3 (N3878, N3874, N2986, N968);
or OR4 (N3879, N3871, N367, N3051, N2910);
buf BUF1 (N3880, N3876);
and AND4 (N3881, N3877, N2153, N587, N1377);
not NOT1 (N3882, N3870);
not NOT1 (N3883, N3882);
not NOT1 (N3884, N3879);
buf BUF1 (N3885, N3880);
and AND2 (N3886, N3883, N167);
not NOT1 (N3887, N3866);
buf BUF1 (N3888, N3885);
nor NOR3 (N3889, N3887, N3624, N1923);
not NOT1 (N3890, N3881);
not NOT1 (N3891, N3884);
nand NAND2 (N3892, N3869, N3575);
nor NOR4 (N3893, N3889, N2880, N3471, N1400);
nand NAND4 (N3894, N3875, N1243, N2611, N1706);
or OR2 (N3895, N3886, N3088);
xor XOR2 (N3896, N3892, N522);
buf BUF1 (N3897, N3878);
nand NAND4 (N3898, N3894, N985, N2482, N934);
nand NAND2 (N3899, N3898, N2261);
nand NAND4 (N3900, N3890, N1669, N1614, N1544);
nor NOR4 (N3901, N3888, N1512, N1121, N2180);
not NOT1 (N3902, N3900);
or OR2 (N3903, N3895, N1690);
not NOT1 (N3904, N3893);
and AND4 (N3905, N3899, N2844, N1345, N2721);
xor XOR2 (N3906, N3896, N3052);
xor XOR2 (N3907, N3891, N1107);
xor XOR2 (N3908, N3873, N2426);
nand NAND4 (N3909, N3903, N1176, N3303, N974);
nor NOR2 (N3910, N3909, N2379);
not NOT1 (N3911, N3901);
buf BUF1 (N3912, N3897);
not NOT1 (N3913, N3911);
not NOT1 (N3914, N3908);
or OR3 (N3915, N3904, N3628, N3492);
buf BUF1 (N3916, N3910);
not NOT1 (N3917, N3913);
nor NOR2 (N3918, N3915, N945);
nand NAND4 (N3919, N3860, N2868, N3052, N511);
buf BUF1 (N3920, N3912);
nor NOR2 (N3921, N3916, N521);
and AND4 (N3922, N3921, N1815, N6, N1527);
or OR3 (N3923, N3906, N20, N2213);
nand NAND2 (N3924, N3902, N3202);
or OR2 (N3925, N3923, N88);
buf BUF1 (N3926, N3914);
or OR4 (N3927, N3926, N3871, N684, N3179);
buf BUF1 (N3928, N3905);
and AND3 (N3929, N3924, N1305, N2910);
not NOT1 (N3930, N3928);
not NOT1 (N3931, N3927);
and AND4 (N3932, N3930, N3097, N3742, N559);
or OR2 (N3933, N3929, N1564);
nand NAND2 (N3934, N3919, N1059);
and AND3 (N3935, N3917, N2720, N900);
or OR3 (N3936, N3932, N3371, N1082);
not NOT1 (N3937, N3935);
xor XOR2 (N3938, N3907, N1188);
xor XOR2 (N3939, N3920, N3089);
nor NOR2 (N3940, N3931, N2174);
nor NOR2 (N3941, N3925, N2966);
nand NAND2 (N3942, N3941, N3677);
nand NAND4 (N3943, N3918, N2134, N3644, N3911);
or OR2 (N3944, N3934, N3376);
not NOT1 (N3945, N3944);
or OR2 (N3946, N3938, N716);
and AND4 (N3947, N3933, N2771, N1094, N1420);
nand NAND3 (N3948, N3947, N2835, N2184);
nor NOR3 (N3949, N3948, N3754, N2111);
nor NOR2 (N3950, N3943, N3151);
not NOT1 (N3951, N3922);
nand NAND3 (N3952, N3950, N1952, N1175);
xor XOR2 (N3953, N3936, N1768);
xor XOR2 (N3954, N3952, N3837);
or OR4 (N3955, N3946, N2508, N3500, N320);
or OR2 (N3956, N3955, N795);
and AND2 (N3957, N3951, N3412);
or OR4 (N3958, N3949, N2556, N1860, N3249);
and AND3 (N3959, N3954, N3016, N2112);
nor NOR2 (N3960, N3937, N1600);
nand NAND3 (N3961, N3940, N1768, N1471);
nand NAND2 (N3962, N3960, N1840);
nor NOR4 (N3963, N3958, N2919, N1961, N3632);
nor NOR3 (N3964, N3942, N3938, N3597);
buf BUF1 (N3965, N3964);
buf BUF1 (N3966, N3962);
not NOT1 (N3967, N3966);
nand NAND2 (N3968, N3939, N2953);
not NOT1 (N3969, N3965);
nand NAND3 (N3970, N3963, N3706, N3136);
xor XOR2 (N3971, N3970, N3766);
nand NAND2 (N3972, N3967, N1113);
not NOT1 (N3973, N3953);
buf BUF1 (N3974, N3969);
and AND3 (N3975, N3971, N3898, N1790);
xor XOR2 (N3976, N3957, N1887);
xor XOR2 (N3977, N3973, N2321);
and AND3 (N3978, N3959, N1201, N2519);
xor XOR2 (N3979, N3945, N2210);
not NOT1 (N3980, N3972);
nor NOR3 (N3981, N3961, N987, N71);
nand NAND2 (N3982, N3975, N3910);
xor XOR2 (N3983, N3977, N619);
nand NAND3 (N3984, N3976, N1981, N3676);
or OR4 (N3985, N3978, N3390, N2901, N858);
and AND3 (N3986, N3983, N2376, N3910);
buf BUF1 (N3987, N3974);
nor NOR2 (N3988, N3979, N1950);
xor XOR2 (N3989, N3982, N1971);
xor XOR2 (N3990, N3988, N1385);
and AND2 (N3991, N3986, N2308);
not NOT1 (N3992, N3987);
xor XOR2 (N3993, N3985, N2510);
nand NAND4 (N3994, N3984, N2383, N363, N3067);
and AND4 (N3995, N3994, N1596, N884, N1052);
buf BUF1 (N3996, N3968);
and AND3 (N3997, N3981, N604, N3036);
nand NAND4 (N3998, N3980, N3129, N1993, N962);
or OR2 (N3999, N3996, N16);
xor XOR2 (N4000, N3998, N2959);
nor NOR4 (N4001, N3997, N2816, N1914, N2948);
nor NOR3 (N4002, N3956, N1321, N2971);
xor XOR2 (N4003, N4000, N2371);
and AND2 (N4004, N3999, N1488);
nor NOR3 (N4005, N4002, N94, N2062);
nor NOR3 (N4006, N3993, N903, N3360);
and AND2 (N4007, N4003, N3376);
buf BUF1 (N4008, N4007);
nor NOR4 (N4009, N4001, N323, N857, N2095);
buf BUF1 (N4010, N3989);
or OR4 (N4011, N4006, N3532, N3857, N2991);
not NOT1 (N4012, N4011);
xor XOR2 (N4013, N3991, N1288);
or OR4 (N4014, N4013, N1258, N578, N2884);
xor XOR2 (N4015, N4004, N406);
nor NOR4 (N4016, N4008, N156, N3686, N2387);
nor NOR2 (N4017, N3992, N2808);
nand NAND2 (N4018, N4010, N1971);
and AND2 (N4019, N4012, N2039);
and AND4 (N4020, N4017, N2449, N689, N3670);
xor XOR2 (N4021, N4015, N3434);
or OR4 (N4022, N4021, N647, N1621, N3154);
not NOT1 (N4023, N4020);
or OR3 (N4024, N4023, N565, N2764);
or OR2 (N4025, N4014, N701);
buf BUF1 (N4026, N4024);
not NOT1 (N4027, N4005);
or OR2 (N4028, N4025, N828);
not NOT1 (N4029, N4016);
nor NOR4 (N4030, N4029, N2575, N3494, N1945);
and AND2 (N4031, N4030, N3653);
nor NOR3 (N4032, N4019, N2180, N2864);
nand NAND4 (N4033, N3990, N271, N762, N1628);
buf BUF1 (N4034, N4033);
xor XOR2 (N4035, N4009, N304);
or OR3 (N4036, N4028, N2460, N677);
and AND2 (N4037, N4031, N1053);
or OR2 (N4038, N3995, N3769);
nor NOR4 (N4039, N4026, N2288, N1032, N736);
nor NOR3 (N4040, N4037, N864, N922);
and AND2 (N4041, N4040, N1289);
xor XOR2 (N4042, N4041, N2602);
and AND3 (N4043, N4018, N472, N2517);
not NOT1 (N4044, N4022);
buf BUF1 (N4045, N4034);
not NOT1 (N4046, N4035);
and AND4 (N4047, N4038, N2787, N2395, N357);
or OR2 (N4048, N4039, N1396);
and AND2 (N4049, N4043, N61);
xor XOR2 (N4050, N4044, N3098);
nand NAND2 (N4051, N4048, N3004);
not NOT1 (N4052, N4046);
and AND3 (N4053, N4042, N3094, N1044);
nand NAND2 (N4054, N4051, N3014);
or OR4 (N4055, N4053, N785, N1561, N3669);
nand NAND2 (N4056, N4055, N2864);
nor NOR3 (N4057, N4054, N4047, N2682);
nand NAND2 (N4058, N1130, N765);
buf BUF1 (N4059, N4032);
and AND4 (N4060, N4049, N2992, N3889, N3217);
nor NOR4 (N4061, N4045, N977, N1579, N3362);
nor NOR4 (N4062, N4050, N442, N4018, N3777);
or OR3 (N4063, N4057, N2498, N1829);
buf BUF1 (N4064, N4059);
not NOT1 (N4065, N4058);
and AND4 (N4066, N4061, N314, N3137, N1858);
xor XOR2 (N4067, N4063, N3731);
nand NAND2 (N4068, N4065, N2594);
and AND3 (N4069, N4068, N2834, N3654);
or OR3 (N4070, N4052, N4029, N1576);
nand NAND2 (N4071, N4062, N2250);
or OR2 (N4072, N4067, N2522);
buf BUF1 (N4073, N4060);
xor XOR2 (N4074, N4066, N2680);
nor NOR3 (N4075, N4069, N1611, N1693);
nand NAND4 (N4076, N4036, N2617, N1586, N398);
or OR4 (N4077, N4070, N1642, N3591, N2020);
not NOT1 (N4078, N4027);
buf BUF1 (N4079, N4056);
and AND2 (N4080, N4073, N697);
nor NOR2 (N4081, N4076, N50);
nand NAND3 (N4082, N4081, N143, N2659);
nand NAND4 (N4083, N4079, N3556, N2752, N2875);
nand NAND3 (N4084, N4083, N1401, N446);
nand NAND2 (N4085, N4074, N1875);
not NOT1 (N4086, N4072);
xor XOR2 (N4087, N4080, N753);
or OR2 (N4088, N4084, N688);
nand NAND4 (N4089, N4086, N1951, N3358, N3546);
nand NAND2 (N4090, N4077, N3824);
and AND4 (N4091, N4088, N1012, N2846, N3353);
nand NAND2 (N4092, N4075, N3609);
and AND4 (N4093, N4092, N3483, N914, N1726);
not NOT1 (N4094, N4090);
nand NAND3 (N4095, N4078, N3833, N3644);
and AND3 (N4096, N4064, N1265, N3650);
buf BUF1 (N4097, N4095);
xor XOR2 (N4098, N4071, N351);
xor XOR2 (N4099, N4085, N2174);
nor NOR2 (N4100, N4082, N2222);
xor XOR2 (N4101, N4089, N376);
not NOT1 (N4102, N4100);
or OR3 (N4103, N4094, N983, N2792);
nand NAND2 (N4104, N4093, N2836);
xor XOR2 (N4105, N4103, N1831);
or OR4 (N4106, N4102, N1724, N2203, N3679);
or OR4 (N4107, N4098, N1143, N2771, N24);
or OR4 (N4108, N4096, N2551, N465, N496);
nand NAND2 (N4109, N4108, N2276);
xor XOR2 (N4110, N4101, N3140);
xor XOR2 (N4111, N4087, N1573);
nor NOR2 (N4112, N4107, N3955);
and AND3 (N4113, N4097, N4041, N2699);
not NOT1 (N4114, N4113);
and AND2 (N4115, N4111, N1298);
nor NOR4 (N4116, N4110, N4107, N1037, N1494);
buf BUF1 (N4117, N4109);
xor XOR2 (N4118, N4099, N1491);
or OR2 (N4119, N4106, N1481);
buf BUF1 (N4120, N4117);
nand NAND4 (N4121, N4115, N191, N2692, N423);
buf BUF1 (N4122, N4112);
buf BUF1 (N4123, N4122);
nor NOR4 (N4124, N4114, N1050, N3499, N11);
xor XOR2 (N4125, N4118, N2188);
not NOT1 (N4126, N4121);
nor NOR2 (N4127, N4105, N2337);
or OR2 (N4128, N4125, N1244);
and AND4 (N4129, N4120, N1024, N3599, N710);
or OR4 (N4130, N4124, N2138, N479, N3495);
and AND3 (N4131, N4129, N3217, N1810);
buf BUF1 (N4132, N4126);
buf BUF1 (N4133, N4116);
nand NAND4 (N4134, N4128, N1373, N866, N1948);
nor NOR4 (N4135, N4127, N3836, N3799, N3419);
xor XOR2 (N4136, N4123, N3562);
buf BUF1 (N4137, N4131);
nor NOR4 (N4138, N4135, N2264, N2836, N151);
nand NAND3 (N4139, N4137, N625, N1886);
nor NOR4 (N4140, N4139, N114, N2407, N3424);
nor NOR4 (N4141, N4130, N56, N2476, N481);
nor NOR3 (N4142, N4119, N2535, N857);
nand NAND2 (N4143, N4136, N2715);
and AND4 (N4144, N4104, N3212, N1925, N2338);
buf BUF1 (N4145, N4143);
or OR3 (N4146, N4145, N1157, N1724);
or OR2 (N4147, N4144, N1462);
buf BUF1 (N4148, N4146);
and AND4 (N4149, N4132, N2013, N51, N3694);
buf BUF1 (N4150, N4149);
and AND4 (N4151, N4150, N3927, N2856, N1402);
buf BUF1 (N4152, N4133);
not NOT1 (N4153, N4140);
and AND4 (N4154, N4152, N3245, N2434, N978);
or OR3 (N4155, N4148, N3372, N1776);
nor NOR3 (N4156, N4153, N2203, N792);
buf BUF1 (N4157, N4155);
nand NAND2 (N4158, N4147, N751);
and AND2 (N4159, N4157, N2586);
nand NAND3 (N4160, N4151, N2222, N1601);
not NOT1 (N4161, N4134);
not NOT1 (N4162, N4091);
nand NAND3 (N4163, N4160, N1664, N2170);
nand NAND4 (N4164, N4162, N770, N3251, N2017);
not NOT1 (N4165, N4158);
nand NAND4 (N4166, N4138, N3134, N4072, N4045);
and AND4 (N4167, N4154, N1618, N953, N1694);
not NOT1 (N4168, N4141);
or OR3 (N4169, N4166, N3764, N138);
nor NOR4 (N4170, N4167, N187, N2781, N2208);
not NOT1 (N4171, N4168);
xor XOR2 (N4172, N4169, N2456);
buf BUF1 (N4173, N4159);
and AND3 (N4174, N4172, N932, N3348);
and AND4 (N4175, N4142, N1869, N475, N2106);
nand NAND3 (N4176, N4170, N2622, N685);
nor NOR4 (N4177, N4161, N3787, N1394, N3926);
nand NAND2 (N4178, N4173, N2392);
or OR2 (N4179, N4177, N2810);
not NOT1 (N4180, N4156);
and AND4 (N4181, N4174, N2223, N4003, N767);
buf BUF1 (N4182, N4171);
and AND3 (N4183, N4179, N2468, N1150);
xor XOR2 (N4184, N4178, N819);
and AND4 (N4185, N4182, N2830, N716, N1728);
and AND3 (N4186, N4180, N3585, N1110);
or OR2 (N4187, N4184, N2124);
not NOT1 (N4188, N4181);
nor NOR3 (N4189, N4185, N48, N232);
nand NAND2 (N4190, N4164, N2257);
buf BUF1 (N4191, N4189);
not NOT1 (N4192, N4163);
not NOT1 (N4193, N4175);
not NOT1 (N4194, N4191);
xor XOR2 (N4195, N4176, N2918);
not NOT1 (N4196, N4195);
nor NOR2 (N4197, N4196, N2096);
and AND3 (N4198, N4194, N891, N3689);
nor NOR4 (N4199, N4183, N1104, N471, N3162);
or OR4 (N4200, N4186, N523, N2437, N2355);
nor NOR2 (N4201, N4192, N3050);
nor NOR2 (N4202, N4165, N601);
and AND3 (N4203, N4201, N4070, N1804);
buf BUF1 (N4204, N4202);
nor NOR3 (N4205, N4203, N2300, N2382);
nor NOR2 (N4206, N4205, N2122);
xor XOR2 (N4207, N4188, N610);
not NOT1 (N4208, N4206);
xor XOR2 (N4209, N4198, N1735);
xor XOR2 (N4210, N4193, N2250);
or OR3 (N4211, N4204, N3033, N240);
buf BUF1 (N4212, N4209);
not NOT1 (N4213, N4187);
and AND3 (N4214, N4207, N489, N2570);
nand NAND4 (N4215, N4212, N2902, N323, N972);
or OR3 (N4216, N4197, N4169, N1274);
or OR2 (N4217, N4199, N2491);
and AND2 (N4218, N4217, N2696);
buf BUF1 (N4219, N4215);
or OR2 (N4220, N4218, N1863);
or OR3 (N4221, N4219, N3221, N3793);
buf BUF1 (N4222, N4190);
not NOT1 (N4223, N4216);
or OR4 (N4224, N4211, N3869, N2695, N3484);
and AND2 (N4225, N4222, N2261);
buf BUF1 (N4226, N4220);
or OR2 (N4227, N4223, N441);
nand NAND3 (N4228, N4210, N2539, N1909);
buf BUF1 (N4229, N4224);
nand NAND4 (N4230, N4214, N2123, N2086, N1688);
nor NOR2 (N4231, N4225, N51);
and AND4 (N4232, N4226, N3956, N2302, N4041);
nand NAND3 (N4233, N4221, N2269, N2315);
buf BUF1 (N4234, N4232);
buf BUF1 (N4235, N4229);
and AND3 (N4236, N4227, N1938, N2484);
not NOT1 (N4237, N4230);
and AND2 (N4238, N4213, N3385);
and AND2 (N4239, N4208, N2549);
nor NOR4 (N4240, N4228, N2440, N3828, N2374);
nand NAND2 (N4241, N4233, N2389);
buf BUF1 (N4242, N4234);
not NOT1 (N4243, N4235);
xor XOR2 (N4244, N4241, N620);
not NOT1 (N4245, N4231);
nor NOR4 (N4246, N4240, N3504, N1496, N599);
or OR3 (N4247, N4246, N3375, N1740);
not NOT1 (N4248, N4247);
or OR2 (N4249, N4200, N250);
xor XOR2 (N4250, N4242, N1437);
and AND2 (N4251, N4243, N3165);
buf BUF1 (N4252, N4237);
and AND3 (N4253, N4249, N1399, N4201);
xor XOR2 (N4254, N4239, N182);
nand NAND2 (N4255, N4238, N2796);
nor NOR2 (N4256, N4236, N2398);
nand NAND3 (N4257, N4256, N3941, N4185);
nor NOR3 (N4258, N4257, N753, N2594);
buf BUF1 (N4259, N4252);
or OR3 (N4260, N4259, N2396, N3947);
or OR3 (N4261, N4248, N2420, N2090);
not NOT1 (N4262, N4260);
nor NOR3 (N4263, N4261, N2548, N958);
buf BUF1 (N4264, N4250);
nand NAND3 (N4265, N4251, N3256, N1670);
xor XOR2 (N4266, N4255, N648);
not NOT1 (N4267, N4264);
nor NOR4 (N4268, N4245, N2255, N1255, N3693);
xor XOR2 (N4269, N4253, N931);
nor NOR3 (N4270, N4262, N1441, N1959);
nand NAND4 (N4271, N4268, N3825, N3609, N2629);
and AND3 (N4272, N4266, N3396, N4124);
or OR2 (N4273, N4267, N922);
xor XOR2 (N4274, N4272, N726);
nand NAND4 (N4275, N4265, N1843, N3524, N2398);
xor XOR2 (N4276, N4254, N4197);
xor XOR2 (N4277, N4269, N2342);
xor XOR2 (N4278, N4277, N3917);
xor XOR2 (N4279, N4274, N2475);
or OR4 (N4280, N4263, N1959, N2661, N1925);
nand NAND4 (N4281, N4276, N281, N65, N3488);
buf BUF1 (N4282, N4281);
and AND2 (N4283, N4271, N849);
xor XOR2 (N4284, N4258, N888);
buf BUF1 (N4285, N4244);
or OR4 (N4286, N4285, N607, N4101, N196);
xor XOR2 (N4287, N4284, N3302);
xor XOR2 (N4288, N4287, N1325);
buf BUF1 (N4289, N4288);
nand NAND2 (N4290, N4280, N1056);
buf BUF1 (N4291, N4278);
and AND4 (N4292, N4282, N3370, N4112, N2769);
buf BUF1 (N4293, N4279);
nor NOR2 (N4294, N4291, N995);
nand NAND2 (N4295, N4294, N1362);
nor NOR2 (N4296, N4273, N725);
not NOT1 (N4297, N4290);
xor XOR2 (N4298, N4297, N698);
buf BUF1 (N4299, N4286);
buf BUF1 (N4300, N4275);
or OR3 (N4301, N4283, N1901, N3024);
buf BUF1 (N4302, N4295);
not NOT1 (N4303, N4296);
and AND2 (N4304, N4292, N2417);
buf BUF1 (N4305, N4303);
and AND4 (N4306, N4298, N3068, N4296, N829);
not NOT1 (N4307, N4305);
nand NAND2 (N4308, N4307, N3164);
or OR4 (N4309, N4293, N2149, N3435, N2133);
not NOT1 (N4310, N4306);
nand NAND4 (N4311, N4270, N1144, N673, N2155);
not NOT1 (N4312, N4309);
buf BUF1 (N4313, N4311);
or OR2 (N4314, N4300, N2032);
buf BUF1 (N4315, N4304);
nor NOR3 (N4316, N4313, N951, N1308);
nand NAND2 (N4317, N4316, N2500);
nand NAND4 (N4318, N4312, N2196, N839, N1387);
nand NAND4 (N4319, N4317, N1636, N1959, N751);
or OR3 (N4320, N4318, N3617, N3207);
not NOT1 (N4321, N4319);
nor NOR3 (N4322, N4299, N4239, N408);
nand NAND3 (N4323, N4301, N2470, N3773);
xor XOR2 (N4324, N4302, N525);
or OR4 (N4325, N4314, N4166, N1243, N2354);
nor NOR3 (N4326, N4322, N1738, N2889);
or OR2 (N4327, N4315, N2898);
not NOT1 (N4328, N4308);
nor NOR4 (N4329, N4324, N4095, N2674, N3241);
and AND2 (N4330, N4325, N828);
xor XOR2 (N4331, N4320, N3824);
not NOT1 (N4332, N4323);
nor NOR4 (N4333, N4289, N2323, N992, N2203);
or OR3 (N4334, N4327, N3869, N2707);
not NOT1 (N4335, N4331);
xor XOR2 (N4336, N4328, N2083);
nor NOR4 (N4337, N4336, N2621, N4163, N1163);
and AND4 (N4338, N4310, N101, N1221, N2326);
buf BUF1 (N4339, N4337);
nor NOR4 (N4340, N4339, N1106, N1651, N4240);
nor NOR2 (N4341, N4332, N4278);
or OR2 (N4342, N4321, N1029);
or OR2 (N4343, N4326, N324);
nor NOR4 (N4344, N4333, N984, N1268, N1642);
xor XOR2 (N4345, N4338, N823);
nand NAND3 (N4346, N4345, N3059, N2159);
xor XOR2 (N4347, N4329, N74);
buf BUF1 (N4348, N4335);
or OR3 (N4349, N4346, N819, N4324);
nand NAND3 (N4350, N4330, N1817, N3146);
nor NOR2 (N4351, N4348, N152);
nor NOR4 (N4352, N4340, N1127, N476, N2210);
nand NAND2 (N4353, N4334, N1953);
buf BUF1 (N4354, N4352);
or OR2 (N4355, N4342, N1392);
buf BUF1 (N4356, N4349);
not NOT1 (N4357, N4350);
and AND2 (N4358, N4343, N4186);
not NOT1 (N4359, N4355);
and AND2 (N4360, N4359, N3550);
nor NOR2 (N4361, N4358, N3203);
not NOT1 (N4362, N4357);
and AND3 (N4363, N4353, N1615, N2463);
or OR2 (N4364, N4344, N1140);
nor NOR4 (N4365, N4361, N3366, N787, N70);
buf BUF1 (N4366, N4365);
not NOT1 (N4367, N4341);
or OR2 (N4368, N4356, N4041);
or OR3 (N4369, N4347, N4116, N982);
nand NAND4 (N4370, N4368, N1166, N4312, N212);
nand NAND3 (N4371, N4369, N1764, N2712);
nor NOR2 (N4372, N4363, N587);
and AND2 (N4373, N4370, N760);
and AND4 (N4374, N4362, N3359, N4099, N674);
and AND2 (N4375, N4354, N3133);
or OR4 (N4376, N4371, N3317, N2224, N1209);
nand NAND4 (N4377, N4373, N1949, N2368, N3078);
nor NOR3 (N4378, N4367, N3243, N1587);
buf BUF1 (N4379, N4376);
nor NOR4 (N4380, N4375, N536, N1438, N1688);
nand NAND4 (N4381, N4366, N3652, N4162, N159);
buf BUF1 (N4382, N4381);
or OR4 (N4383, N4364, N1899, N3107, N2783);
nor NOR3 (N4384, N4374, N2859, N1830);
nand NAND2 (N4385, N4379, N2591);
buf BUF1 (N4386, N4383);
or OR4 (N4387, N4385, N4091, N2636, N3347);
and AND4 (N4388, N4351, N499, N1922, N388);
nor NOR3 (N4389, N4387, N2826, N2450);
and AND3 (N4390, N4386, N1666, N2803);
buf BUF1 (N4391, N4378);
and AND4 (N4392, N4372, N2603, N3903, N3961);
and AND4 (N4393, N4384, N624, N841, N115);
not NOT1 (N4394, N4380);
nor NOR4 (N4395, N4393, N491, N3365, N4360);
buf BUF1 (N4396, N1289);
and AND2 (N4397, N4395, N488);
or OR2 (N4398, N4388, N278);
nor NOR3 (N4399, N4382, N4043, N1092);
xor XOR2 (N4400, N4392, N3266);
and AND2 (N4401, N4397, N837);
not NOT1 (N4402, N4390);
xor XOR2 (N4403, N4400, N4022);
nor NOR4 (N4404, N4394, N3828, N1603, N66);
not NOT1 (N4405, N4398);
and AND3 (N4406, N4402, N170, N406);
and AND4 (N4407, N4403, N844, N3556, N3300);
and AND2 (N4408, N4377, N1355);
nor NOR3 (N4409, N4408, N159, N1059);
buf BUF1 (N4410, N4407);
or OR3 (N4411, N4409, N2835, N1038);
xor XOR2 (N4412, N4401, N3067);
not NOT1 (N4413, N4389);
or OR3 (N4414, N4405, N1833, N4364);
nand NAND4 (N4415, N4399, N459, N3777, N3791);
and AND4 (N4416, N4412, N1302, N3353, N3329);
buf BUF1 (N4417, N4406);
nor NOR3 (N4418, N4414, N669, N2184);
buf BUF1 (N4419, N4411);
not NOT1 (N4420, N4391);
nor NOR4 (N4421, N4418, N703, N2921, N2420);
nand NAND4 (N4422, N4419, N645, N337, N3510);
xor XOR2 (N4423, N4421, N1394);
nor NOR3 (N4424, N4423, N1211, N2887);
or OR2 (N4425, N4422, N2380);
buf BUF1 (N4426, N4417);
not NOT1 (N4427, N4415);
or OR2 (N4428, N4404, N1222);
and AND2 (N4429, N4396, N2125);
xor XOR2 (N4430, N4429, N1513);
or OR2 (N4431, N4427, N3717);
nand NAND2 (N4432, N4410, N3189);
or OR3 (N4433, N4420, N1187, N354);
buf BUF1 (N4434, N4428);
xor XOR2 (N4435, N4425, N1298);
nor NOR3 (N4436, N4424, N3357, N3333);
or OR2 (N4437, N4432, N2440);
buf BUF1 (N4438, N4434);
nand NAND4 (N4439, N4437, N4393, N3238, N786);
nor NOR2 (N4440, N4436, N3043);
not NOT1 (N4441, N4435);
nand NAND3 (N4442, N4426, N4087, N2538);
buf BUF1 (N4443, N4431);
and AND4 (N4444, N4440, N2586, N2348, N2480);
not NOT1 (N4445, N4430);
nand NAND2 (N4446, N4416, N3638);
nand NAND3 (N4447, N4433, N2894, N3583);
or OR2 (N4448, N4445, N244);
nor NOR3 (N4449, N4447, N974, N3180);
or OR2 (N4450, N4444, N4079);
not NOT1 (N4451, N4441);
buf BUF1 (N4452, N4413);
and AND2 (N4453, N4449, N1103);
and AND3 (N4454, N4450, N1646, N2930);
nor NOR3 (N4455, N4452, N1957, N1996);
nor NOR2 (N4456, N4451, N1667);
buf BUF1 (N4457, N4443);
and AND2 (N4458, N4456, N197);
not NOT1 (N4459, N4458);
not NOT1 (N4460, N4438);
xor XOR2 (N4461, N4446, N3628);
nor NOR2 (N4462, N4439, N489);
nand NAND4 (N4463, N4454, N4094, N1785, N287);
and AND4 (N4464, N4442, N4258, N3978, N825);
or OR2 (N4465, N4457, N3652);
xor XOR2 (N4466, N4461, N2754);
or OR3 (N4467, N4466, N2511, N3253);
and AND2 (N4468, N4460, N4348);
or OR2 (N4469, N4465, N3130);
or OR2 (N4470, N4464, N4154);
or OR4 (N4471, N4462, N2617, N4421, N839);
and AND3 (N4472, N4459, N1574, N1725);
or OR3 (N4473, N4470, N3737, N3907);
nand NAND2 (N4474, N4468, N3550);
nand NAND2 (N4475, N4463, N1490);
xor XOR2 (N4476, N4471, N4313);
nand NAND4 (N4477, N4469, N4435, N1226, N4059);
nand NAND4 (N4478, N4473, N1392, N40, N4180);
nand NAND4 (N4479, N4453, N3107, N1483, N1381);
and AND2 (N4480, N4455, N1843);
not NOT1 (N4481, N4477);
and AND4 (N4482, N4478, N881, N329, N1241);
nand NAND4 (N4483, N4474, N2740, N4069, N4051);
or OR4 (N4484, N4475, N1514, N315, N208);
nand NAND4 (N4485, N4479, N3651, N1178, N1553);
xor XOR2 (N4486, N4480, N1944);
xor XOR2 (N4487, N4476, N1671);
and AND4 (N4488, N4486, N2408, N4113, N3267);
or OR3 (N4489, N4487, N1474, N4060);
and AND4 (N4490, N4489, N1601, N1356, N982);
not NOT1 (N4491, N4482);
xor XOR2 (N4492, N4485, N2830);
nand NAND3 (N4493, N4484, N1883, N1891);
not NOT1 (N4494, N4448);
nor NOR3 (N4495, N4493, N1655, N3267);
and AND4 (N4496, N4492, N2462, N2702, N1560);
and AND4 (N4497, N4481, N3204, N1087, N4452);
or OR4 (N4498, N4472, N2763, N3665, N1711);
or OR2 (N4499, N4488, N4265);
and AND3 (N4500, N4467, N2953, N4469);
or OR4 (N4501, N4496, N1337, N1049, N1943);
or OR4 (N4502, N4501, N927, N1073, N3889);
not NOT1 (N4503, N4494);
xor XOR2 (N4504, N4495, N3800);
or OR4 (N4505, N4500, N4454, N1954, N443);
or OR2 (N4506, N4491, N4158);
buf BUF1 (N4507, N4499);
and AND3 (N4508, N4502, N4434, N401);
not NOT1 (N4509, N4498);
or OR3 (N4510, N4497, N1035, N3845);
nand NAND4 (N4511, N4508, N3329, N405, N3165);
nand NAND4 (N4512, N4503, N1135, N4075, N2859);
xor XOR2 (N4513, N4509, N1359);
or OR2 (N4514, N4512, N4356);
buf BUF1 (N4515, N4511);
or OR3 (N4516, N4506, N655, N2566);
not NOT1 (N4517, N4505);
xor XOR2 (N4518, N4504, N612);
not NOT1 (N4519, N4517);
buf BUF1 (N4520, N4518);
buf BUF1 (N4521, N4520);
or OR2 (N4522, N4483, N3509);
nand NAND2 (N4523, N4521, N4093);
or OR4 (N4524, N4519, N3216, N2706, N4258);
buf BUF1 (N4525, N4515);
buf BUF1 (N4526, N4522);
and AND3 (N4527, N4523, N1428, N644);
xor XOR2 (N4528, N4514, N47);
or OR2 (N4529, N4524, N1526);
nand NAND4 (N4530, N4527, N2881, N855, N608);
nor NOR2 (N4531, N4528, N3119);
nor NOR3 (N4532, N4507, N3708, N1287);
and AND4 (N4533, N4531, N4397, N2046, N3117);
buf BUF1 (N4534, N4513);
not NOT1 (N4535, N4490);
not NOT1 (N4536, N4525);
nand NAND4 (N4537, N4529, N1884, N2467, N2505);
nand NAND2 (N4538, N4533, N1154);
and AND2 (N4539, N4526, N41);
buf BUF1 (N4540, N4536);
xor XOR2 (N4541, N4530, N2601);
buf BUF1 (N4542, N4516);
nor NOR3 (N4543, N4539, N2132, N220);
nand NAND4 (N4544, N4543, N2599, N1260, N3049);
xor XOR2 (N4545, N4537, N788);
nand NAND4 (N4546, N4544, N2578, N2407, N3872);
or OR3 (N4547, N4540, N2074, N3942);
not NOT1 (N4548, N4542);
nor NOR4 (N4549, N4546, N4261, N4222, N62);
nor NOR4 (N4550, N4548, N2013, N3406, N1302);
not NOT1 (N4551, N4541);
buf BUF1 (N4552, N4545);
nand NAND2 (N4553, N4532, N4230);
nand NAND2 (N4554, N4552, N3);
and AND3 (N4555, N4554, N3028, N3372);
buf BUF1 (N4556, N4553);
buf BUF1 (N4557, N4555);
not NOT1 (N4558, N4535);
buf BUF1 (N4559, N4551);
nand NAND4 (N4560, N4550, N2393, N942, N3039);
not NOT1 (N4561, N4556);
not NOT1 (N4562, N4559);
not NOT1 (N4563, N4562);
nor NOR4 (N4564, N4549, N939, N3348, N3165);
nand NAND2 (N4565, N4558, N73);
and AND4 (N4566, N4564, N3218, N177, N788);
nor NOR4 (N4567, N4565, N3452, N1532, N2159);
not NOT1 (N4568, N4560);
nand NAND4 (N4569, N4547, N661, N173, N2597);
nand NAND4 (N4570, N4566, N3653, N270, N2981);
and AND3 (N4571, N4510, N3834, N311);
or OR2 (N4572, N4568, N256);
buf BUF1 (N4573, N4534);
and AND2 (N4574, N4563, N3079);
nand NAND2 (N4575, N4538, N751);
not NOT1 (N4576, N4575);
or OR2 (N4577, N4567, N1330);
nor NOR3 (N4578, N4577, N601, N1143);
or OR4 (N4579, N4569, N2950, N2284, N721);
nand NAND4 (N4580, N4576, N3266, N4078, N3324);
and AND4 (N4581, N4579, N2604, N753, N2815);
xor XOR2 (N4582, N4573, N3572);
nor NOR4 (N4583, N4581, N3437, N4477, N1296);
nand NAND3 (N4584, N4557, N4382, N1636);
nor NOR3 (N4585, N4582, N438, N4490);
or OR4 (N4586, N4585, N2938, N2809, N1542);
buf BUF1 (N4587, N4584);
buf BUF1 (N4588, N4583);
not NOT1 (N4589, N4580);
not NOT1 (N4590, N4561);
nor NOR2 (N4591, N4574, N2157);
xor XOR2 (N4592, N4590, N2464);
nand NAND3 (N4593, N4578, N545, N1192);
buf BUF1 (N4594, N4571);
nand NAND4 (N4595, N4587, N26, N63, N4363);
nand NAND2 (N4596, N4594, N2110);
not NOT1 (N4597, N4589);
and AND3 (N4598, N4572, N3203, N2659);
xor XOR2 (N4599, N4586, N2046);
and AND2 (N4600, N4570, N592);
and AND3 (N4601, N4591, N307, N4215);
nand NAND3 (N4602, N4593, N1870, N3387);
nand NAND4 (N4603, N4600, N576, N2552, N3426);
and AND4 (N4604, N4595, N2166, N899, N2693);
not NOT1 (N4605, N4599);
buf BUF1 (N4606, N4597);
not NOT1 (N4607, N4602);
and AND3 (N4608, N4596, N2916, N4463);
not NOT1 (N4609, N4604);
not NOT1 (N4610, N4601);
or OR4 (N4611, N4609, N3011, N3203, N2553);
xor XOR2 (N4612, N4610, N1747);
nor NOR4 (N4613, N4588, N784, N3254, N3858);
or OR4 (N4614, N4598, N3094, N3118, N646);
nor NOR3 (N4615, N4592, N737, N1169);
buf BUF1 (N4616, N4603);
not NOT1 (N4617, N4611);
not NOT1 (N4618, N4616);
not NOT1 (N4619, N4612);
not NOT1 (N4620, N4607);
not NOT1 (N4621, N4619);
xor XOR2 (N4622, N4621, N3683);
or OR2 (N4623, N4608, N408);
and AND4 (N4624, N4605, N4075, N400, N4089);
not NOT1 (N4625, N4622);
nand NAND2 (N4626, N4625, N3661);
not NOT1 (N4627, N4606);
xor XOR2 (N4628, N4617, N2306);
nand NAND3 (N4629, N4627, N2112, N246);
xor XOR2 (N4630, N4620, N2181);
buf BUF1 (N4631, N4615);
nand NAND4 (N4632, N4629, N233, N1659, N3227);
not NOT1 (N4633, N4618);
buf BUF1 (N4634, N4631);
or OR3 (N4635, N4628, N1269, N2685);
and AND3 (N4636, N4614, N2527, N4620);
not NOT1 (N4637, N4630);
nand NAND4 (N4638, N4626, N2775, N1676, N1728);
xor XOR2 (N4639, N4633, N4365);
nand NAND4 (N4640, N4638, N101, N1165, N623);
and AND3 (N4641, N4634, N2742, N3163);
or OR4 (N4642, N4624, N3410, N1912, N1258);
or OR3 (N4643, N4639, N119, N1205);
or OR3 (N4644, N4636, N4452, N1683);
or OR3 (N4645, N4613, N710, N374);
or OR2 (N4646, N4640, N2860);
xor XOR2 (N4647, N4646, N3779);
xor XOR2 (N4648, N4641, N732);
and AND2 (N4649, N4645, N2629);
not NOT1 (N4650, N4643);
xor XOR2 (N4651, N4632, N246);
buf BUF1 (N4652, N4623);
not NOT1 (N4653, N4650);
not NOT1 (N4654, N4642);
xor XOR2 (N4655, N4654, N2095);
xor XOR2 (N4656, N4648, N835);
and AND2 (N4657, N4635, N3302);
not NOT1 (N4658, N4652);
and AND4 (N4659, N4656, N679, N2329, N3792);
or OR2 (N4660, N4644, N2019);
not NOT1 (N4661, N4660);
xor XOR2 (N4662, N4659, N3575);
xor XOR2 (N4663, N4653, N4394);
nand NAND2 (N4664, N4655, N3652);
nor NOR2 (N4665, N4664, N822);
nand NAND2 (N4666, N4657, N2600);
not NOT1 (N4667, N4658);
not NOT1 (N4668, N4637);
nor NOR3 (N4669, N4663, N2995, N2058);
or OR3 (N4670, N4667, N3682, N2418);
or OR4 (N4671, N4662, N1470, N1610, N127);
not NOT1 (N4672, N4647);
not NOT1 (N4673, N4669);
nor NOR2 (N4674, N4661, N2497);
or OR3 (N4675, N4666, N494, N892);
nand NAND4 (N4676, N4668, N4508, N1724, N349);
not NOT1 (N4677, N4665);
xor XOR2 (N4678, N4651, N1523);
xor XOR2 (N4679, N4677, N4465);
xor XOR2 (N4680, N4675, N3);
and AND4 (N4681, N4670, N1700, N4171, N2654);
and AND4 (N4682, N4671, N1504, N3134, N3793);
nor NOR2 (N4683, N4674, N3663);
or OR2 (N4684, N4672, N3743);
nand NAND3 (N4685, N4681, N3408, N103);
nor NOR4 (N4686, N4680, N2165, N2820, N4334);
or OR4 (N4687, N4682, N2275, N496, N4207);
buf BUF1 (N4688, N4686);
xor XOR2 (N4689, N4683, N649);
nand NAND2 (N4690, N4679, N3167);
and AND2 (N4691, N4649, N988);
not NOT1 (N4692, N4690);
xor XOR2 (N4693, N4689, N2249);
or OR3 (N4694, N4684, N3733, N66);
and AND4 (N4695, N4688, N878, N4399, N1725);
xor XOR2 (N4696, N4676, N373);
nand NAND4 (N4697, N4695, N1478, N4400, N220);
buf BUF1 (N4698, N4696);
nand NAND4 (N4699, N4673, N2726, N328, N2058);
not NOT1 (N4700, N4692);
not NOT1 (N4701, N4678);
and AND4 (N4702, N4700, N3533, N2960, N1093);
nor NOR2 (N4703, N4685, N83);
xor XOR2 (N4704, N4691, N4497);
nand NAND4 (N4705, N4693, N598, N1029, N1076);
or OR4 (N4706, N4702, N96, N2436, N1645);
and AND4 (N4707, N4705, N1609, N24, N4614);
xor XOR2 (N4708, N4687, N2415);
buf BUF1 (N4709, N4699);
nand NAND3 (N4710, N4694, N1090, N4163);
nor NOR2 (N4711, N4697, N3994);
buf BUF1 (N4712, N4709);
buf BUF1 (N4713, N4704);
buf BUF1 (N4714, N4711);
xor XOR2 (N4715, N4714, N1820);
xor XOR2 (N4716, N4712, N1437);
or OR2 (N4717, N4701, N3807);
xor XOR2 (N4718, N4707, N2459);
nand NAND2 (N4719, N4703, N1510);
or OR2 (N4720, N4715, N3256);
buf BUF1 (N4721, N4718);
nor NOR3 (N4722, N4716, N2560, N2682);
nand NAND3 (N4723, N4713, N2566, N2115);
xor XOR2 (N4724, N4710, N2242);
xor XOR2 (N4725, N4720, N2535);
nor NOR2 (N4726, N4698, N118);
nand NAND2 (N4727, N4721, N145);
not NOT1 (N4728, N4717);
or OR2 (N4729, N4722, N1120);
or OR4 (N4730, N4719, N2007, N3767, N3698);
or OR4 (N4731, N4726, N3883, N1793, N4159);
and AND3 (N4732, N4729, N4595, N3449);
nor NOR3 (N4733, N4725, N1019, N598);
buf BUF1 (N4734, N4708);
and AND4 (N4735, N4724, N4351, N906, N4543);
not NOT1 (N4736, N4727);
and AND4 (N4737, N4728, N4365, N243, N568);
xor XOR2 (N4738, N4737, N2988);
and AND3 (N4739, N4723, N1346, N1195);
buf BUF1 (N4740, N4734);
xor XOR2 (N4741, N4735, N1441);
nor NOR3 (N4742, N4731, N650, N3154);
buf BUF1 (N4743, N4706);
not NOT1 (N4744, N4740);
xor XOR2 (N4745, N4744, N1855);
nor NOR4 (N4746, N4738, N3474, N1378, N34);
nor NOR4 (N4747, N4743, N1899, N1083, N3944);
xor XOR2 (N4748, N4739, N285);
or OR2 (N4749, N4748, N73);
nand NAND2 (N4750, N4741, N3884);
xor XOR2 (N4751, N4742, N2022);
and AND3 (N4752, N4730, N2590, N4138);
nand NAND4 (N4753, N4747, N662, N2923, N69);
xor XOR2 (N4754, N4736, N2137);
xor XOR2 (N4755, N4732, N2682);
nand NAND3 (N4756, N4753, N665, N1317);
nor NOR2 (N4757, N4745, N2349);
xor XOR2 (N4758, N4755, N1757);
xor XOR2 (N4759, N4756, N4622);
xor XOR2 (N4760, N4749, N3596);
and AND3 (N4761, N4758, N1901, N4172);
and AND4 (N4762, N4754, N2438, N4735, N1643);
and AND3 (N4763, N4761, N1908, N4496);
nand NAND3 (N4764, N4757, N3096, N2161);
and AND2 (N4765, N4752, N1245);
nand NAND2 (N4766, N4760, N4461);
buf BUF1 (N4767, N4764);
and AND3 (N4768, N4765, N3302, N3699);
nor NOR4 (N4769, N4751, N626, N3149, N4334);
or OR2 (N4770, N4769, N3253);
xor XOR2 (N4771, N4733, N3868);
not NOT1 (N4772, N4759);
xor XOR2 (N4773, N4766, N317);
or OR3 (N4774, N4762, N4521, N864);
buf BUF1 (N4775, N4763);
nand NAND4 (N4776, N4774, N964, N1187, N830);
buf BUF1 (N4777, N4772);
not NOT1 (N4778, N4776);
xor XOR2 (N4779, N4768, N449);
or OR4 (N4780, N4770, N2843, N2388, N1287);
buf BUF1 (N4781, N4779);
buf BUF1 (N4782, N4771);
nor NOR2 (N4783, N4781, N4031);
xor XOR2 (N4784, N4780, N3428);
and AND3 (N4785, N4782, N497, N399);
nor NOR2 (N4786, N4785, N986);
or OR3 (N4787, N4783, N1974, N1996);
nand NAND2 (N4788, N4773, N1902);
xor XOR2 (N4789, N4788, N4165);
nand NAND3 (N4790, N4786, N301, N1749);
not NOT1 (N4791, N4789);
and AND2 (N4792, N4775, N614);
xor XOR2 (N4793, N4791, N307);
nor NOR3 (N4794, N4790, N203, N744);
buf BUF1 (N4795, N4794);
not NOT1 (N4796, N4750);
or OR2 (N4797, N4787, N785);
not NOT1 (N4798, N4746);
nand NAND4 (N4799, N4778, N169, N116, N1268);
nor NOR3 (N4800, N4799, N4755, N650);
buf BUF1 (N4801, N4777);
not NOT1 (N4802, N4798);
buf BUF1 (N4803, N4784);
nor NOR2 (N4804, N4802, N4052);
xor XOR2 (N4805, N4801, N4545);
xor XOR2 (N4806, N4803, N2082);
or OR4 (N4807, N4797, N602, N4366, N643);
and AND3 (N4808, N4795, N2265, N1080);
buf BUF1 (N4809, N4804);
not NOT1 (N4810, N4800);
nor NOR2 (N4811, N4808, N1287);
not NOT1 (N4812, N4811);
nor NOR3 (N4813, N4806, N3338, N1514);
buf BUF1 (N4814, N4793);
or OR4 (N4815, N4810, N4014, N2410, N1011);
nand NAND4 (N4816, N4813, N4743, N1492, N72);
nor NOR4 (N4817, N4812, N2080, N4325, N3657);
and AND2 (N4818, N4817, N4437);
and AND2 (N4819, N4815, N4041);
and AND4 (N4820, N4805, N3194, N1169, N3595);
or OR4 (N4821, N4818, N503, N4198, N2491);
nand NAND4 (N4822, N4821, N3581, N1840, N2624);
xor XOR2 (N4823, N4809, N3400);
or OR4 (N4824, N4792, N4427, N3183, N2557);
not NOT1 (N4825, N4819);
not NOT1 (N4826, N4767);
not NOT1 (N4827, N4823);
and AND4 (N4828, N4825, N3169, N1742, N1798);
buf BUF1 (N4829, N4826);
not NOT1 (N4830, N4822);
not NOT1 (N4831, N4820);
buf BUF1 (N4832, N4827);
nor NOR4 (N4833, N4816, N2898, N2959, N71);
or OR2 (N4834, N4807, N161);
and AND3 (N4835, N4814, N3746, N4248);
xor XOR2 (N4836, N4828, N4646);
xor XOR2 (N4837, N4835, N4212);
nor NOR3 (N4838, N4796, N4704, N399);
xor XOR2 (N4839, N4831, N2148);
not NOT1 (N4840, N4833);
buf BUF1 (N4841, N4836);
or OR4 (N4842, N4837, N2556, N3796, N2372);
or OR4 (N4843, N4824, N3127, N2590, N3370);
not NOT1 (N4844, N4838);
and AND2 (N4845, N4842, N2262);
not NOT1 (N4846, N4832);
nand NAND3 (N4847, N4844, N980, N1894);
buf BUF1 (N4848, N4847);
not NOT1 (N4849, N4834);
or OR3 (N4850, N4840, N1794, N2946);
nor NOR3 (N4851, N4829, N2152, N2517);
or OR2 (N4852, N4846, N3463);
or OR4 (N4853, N4830, N594, N1913, N1859);
or OR2 (N4854, N4850, N3561);
nor NOR3 (N4855, N4843, N1630, N170);
nand NAND2 (N4856, N4841, N4057);
nor NOR2 (N4857, N4852, N1213);
and AND4 (N4858, N4856, N4668, N3193, N761);
and AND3 (N4859, N4849, N1510, N1262);
not NOT1 (N4860, N4848);
xor XOR2 (N4861, N4845, N4295);
or OR3 (N4862, N4853, N1999, N660);
nor NOR2 (N4863, N4861, N4565);
nor NOR4 (N4864, N4858, N1691, N6, N3407);
buf BUF1 (N4865, N4864);
not NOT1 (N4866, N4862);
or OR4 (N4867, N4854, N608, N125, N59);
xor XOR2 (N4868, N4866, N906);
xor XOR2 (N4869, N4839, N4544);
not NOT1 (N4870, N4869);
or OR4 (N4871, N4865, N898, N3484, N856);
or OR4 (N4872, N4859, N2362, N2721, N1058);
or OR2 (N4873, N4857, N2733);
and AND3 (N4874, N4873, N1680, N1725);
or OR4 (N4875, N4855, N1489, N1070, N3256);
or OR2 (N4876, N4871, N3590);
not NOT1 (N4877, N4863);
not NOT1 (N4878, N4877);
xor XOR2 (N4879, N4851, N1461);
nand NAND4 (N4880, N4879, N4533, N331, N114);
or OR3 (N4881, N4880, N3000, N859);
and AND3 (N4882, N4875, N3399, N2979);
and AND2 (N4883, N4882, N1258);
or OR4 (N4884, N4874, N471, N3884, N3489);
nor NOR4 (N4885, N4868, N1117, N1513, N3395);
xor XOR2 (N4886, N4884, N3544);
xor XOR2 (N4887, N4876, N574);
and AND3 (N4888, N4867, N3296, N1690);
buf BUF1 (N4889, N4860);
nand NAND3 (N4890, N4872, N3727, N4770);
and AND3 (N4891, N4890, N1325, N607);
nor NOR4 (N4892, N4886, N2810, N4249, N1480);
not NOT1 (N4893, N4888);
and AND4 (N4894, N4892, N3594, N4306, N3021);
nand NAND3 (N4895, N4870, N4609, N210);
nand NAND4 (N4896, N4889, N2537, N4080, N2223);
not NOT1 (N4897, N4893);
or OR3 (N4898, N4897, N3394, N2815);
not NOT1 (N4899, N4878);
buf BUF1 (N4900, N4896);
nand NAND3 (N4901, N4883, N2299, N772);
buf BUF1 (N4902, N4885);
nor NOR3 (N4903, N4902, N2962, N1026);
not NOT1 (N4904, N4898);
and AND3 (N4905, N4899, N291, N1637);
not NOT1 (N4906, N4895);
or OR3 (N4907, N4881, N1729, N4654);
not NOT1 (N4908, N4906);
nor NOR3 (N4909, N4901, N2762, N2274);
buf BUF1 (N4910, N4908);
not NOT1 (N4911, N4905);
nor NOR2 (N4912, N4907, N4371);
and AND4 (N4913, N4912, N3932, N408, N3983);
buf BUF1 (N4914, N4913);
nor NOR4 (N4915, N4904, N1422, N2399, N3546);
and AND2 (N4916, N4911, N3270);
nor NOR4 (N4917, N4894, N753, N1618, N2733);
buf BUF1 (N4918, N4900);
not NOT1 (N4919, N4917);
nand NAND4 (N4920, N4887, N3360, N1806, N1558);
buf BUF1 (N4921, N4915);
nor NOR2 (N4922, N4920, N2591);
not NOT1 (N4923, N4909);
buf BUF1 (N4924, N4921);
and AND4 (N4925, N4903, N177, N3657, N130);
and AND3 (N4926, N4891, N376, N2767);
or OR3 (N4927, N4916, N2626, N3635);
or OR4 (N4928, N4926, N3631, N408, N1146);
nand NAND2 (N4929, N4924, N3453);
xor XOR2 (N4930, N4914, N2275);
xor XOR2 (N4931, N4925, N777);
buf BUF1 (N4932, N4928);
nor NOR4 (N4933, N4927, N1107, N1131, N3034);
nor NOR4 (N4934, N4930, N4280, N4239, N3246);
not NOT1 (N4935, N4918);
xor XOR2 (N4936, N4923, N287);
not NOT1 (N4937, N4935);
or OR4 (N4938, N4936, N661, N4256, N3534);
buf BUF1 (N4939, N4929);
nand NAND2 (N4940, N4922, N2297);
nand NAND2 (N4941, N4919, N2949);
nand NAND2 (N4942, N4939, N2263);
and AND3 (N4943, N4938, N3904, N589);
xor XOR2 (N4944, N4937, N171);
buf BUF1 (N4945, N4940);
and AND4 (N4946, N4931, N248, N3313, N4709);
buf BUF1 (N4947, N4946);
or OR2 (N4948, N4942, N1835);
nor NOR4 (N4949, N4945, N397, N2457, N4512);
nand NAND3 (N4950, N4944, N309, N3581);
buf BUF1 (N4951, N4934);
xor XOR2 (N4952, N4947, N2628);
not NOT1 (N4953, N4948);
nor NOR3 (N4954, N4943, N275, N330);
nor NOR3 (N4955, N4910, N150, N2348);
or OR3 (N4956, N4952, N733, N2494);
xor XOR2 (N4957, N4932, N4691);
not NOT1 (N4958, N4949);
or OR2 (N4959, N4954, N1808);
buf BUF1 (N4960, N4958);
nor NOR4 (N4961, N4957, N2820, N3192, N732);
nor NOR2 (N4962, N4959, N4248);
and AND2 (N4963, N4955, N2174);
or OR3 (N4964, N4963, N514, N3293);
buf BUF1 (N4965, N4961);
nand NAND4 (N4966, N4960, N212, N1175, N2335);
nor NOR3 (N4967, N4953, N3428, N743);
buf BUF1 (N4968, N4966);
xor XOR2 (N4969, N4965, N2619);
nand NAND4 (N4970, N4967, N4370, N1859, N3077);
and AND2 (N4971, N4962, N1253);
buf BUF1 (N4972, N4941);
and AND3 (N4973, N4956, N94, N3875);
buf BUF1 (N4974, N4973);
not NOT1 (N4975, N4970);
nand NAND4 (N4976, N4933, N4358, N3175, N3556);
or OR4 (N4977, N4976, N321, N4717, N3366);
or OR2 (N4978, N4977, N4516);
or OR3 (N4979, N4978, N4291, N3174);
or OR3 (N4980, N4972, N3202, N3931);
and AND3 (N4981, N4975, N2565, N1486);
and AND2 (N4982, N4950, N4879);
or OR2 (N4983, N4974, N2916);
xor XOR2 (N4984, N4964, N768);
and AND4 (N4985, N4971, N760, N765, N1726);
buf BUF1 (N4986, N4984);
nor NOR4 (N4987, N4985, N191, N2613, N4050);
nor NOR2 (N4988, N4980, N2736);
or OR4 (N4989, N4988, N3210, N4430, N4924);
not NOT1 (N4990, N4982);
and AND4 (N4991, N4987, N2599, N1381, N2080);
xor XOR2 (N4992, N4979, N4854);
xor XOR2 (N4993, N4991, N4093);
not NOT1 (N4994, N4969);
nand NAND2 (N4995, N4951, N262);
xor XOR2 (N4996, N4992, N3680);
nand NAND3 (N4997, N4994, N1153, N475);
not NOT1 (N4998, N4983);
xor XOR2 (N4999, N4998, N850);
nand NAND2 (N5000, N4989, N3389);
nor NOR2 (N5001, N5000, N4325);
nand NAND3 (N5002, N5001, N1890, N4641);
or OR2 (N5003, N4993, N4481);
or OR4 (N5004, N4986, N1210, N3934, N496);
not NOT1 (N5005, N4968);
buf BUF1 (N5006, N4995);
not NOT1 (N5007, N5002);
nand NAND4 (N5008, N4997, N3854, N1675, N748);
or OR4 (N5009, N5007, N3083, N4207, N961);
buf BUF1 (N5010, N5005);
not NOT1 (N5011, N5004);
and AND3 (N5012, N5008, N3787, N1811);
not NOT1 (N5013, N4999);
buf BUF1 (N5014, N5013);
and AND3 (N5015, N5012, N1487, N3685);
or OR4 (N5016, N5010, N4459, N2534, N1330);
nor NOR2 (N5017, N4990, N18);
nand NAND2 (N5018, N5009, N1549);
and AND3 (N5019, N5018, N3468, N3712);
and AND4 (N5020, N4981, N846, N1278, N4713);
buf BUF1 (N5021, N5011);
and AND2 (N5022, N5017, N3962);
not NOT1 (N5023, N5016);
nor NOR4 (N5024, N5003, N490, N3593, N3635);
not NOT1 (N5025, N5020);
nand NAND4 (N5026, N5024, N2333, N1490, N4053);
or OR3 (N5027, N5025, N2039, N1501);
not NOT1 (N5028, N5021);
nor NOR3 (N5029, N5019, N2815, N1251);
nand NAND4 (N5030, N5027, N713, N525, N794);
and AND2 (N5031, N5028, N1644);
nand NAND3 (N5032, N5030, N490, N264);
xor XOR2 (N5033, N5031, N3025);
buf BUF1 (N5034, N5033);
xor XOR2 (N5035, N5023, N4950);
and AND4 (N5036, N5014, N3131, N4968, N3143);
or OR2 (N5037, N5032, N1164);
xor XOR2 (N5038, N5037, N1916);
not NOT1 (N5039, N5038);
and AND2 (N5040, N5015, N4565);
not NOT1 (N5041, N5029);
xor XOR2 (N5042, N5034, N1959);
nor NOR4 (N5043, N4996, N4816, N443, N1504);
xor XOR2 (N5044, N5006, N2553);
xor XOR2 (N5045, N5040, N79);
not NOT1 (N5046, N5035);
buf BUF1 (N5047, N5045);
nor NOR4 (N5048, N5036, N4024, N182, N626);
xor XOR2 (N5049, N5041, N3976);
xor XOR2 (N5050, N5026, N3144);
and AND2 (N5051, N5047, N2318);
buf BUF1 (N5052, N5022);
nor NOR3 (N5053, N5043, N2000, N478);
nand NAND3 (N5054, N5052, N3895, N3928);
nor NOR2 (N5055, N5050, N1197);
nand NAND4 (N5056, N5049, N1774, N773, N3620);
not NOT1 (N5057, N5039);
and AND4 (N5058, N5056, N3599, N554, N777);
nor NOR2 (N5059, N5051, N240);
nand NAND4 (N5060, N5042, N1646, N4277, N3849);
buf BUF1 (N5061, N5055);
nor NOR4 (N5062, N5061, N4064, N1969, N4968);
not NOT1 (N5063, N5048);
and AND4 (N5064, N5058, N1162, N4863, N2029);
or OR4 (N5065, N5062, N4931, N2031, N2680);
or OR3 (N5066, N5046, N4148, N3189);
or OR3 (N5067, N5064, N1132, N4387);
or OR2 (N5068, N5060, N2501);
and AND4 (N5069, N5059, N3614, N484, N250);
xor XOR2 (N5070, N5057, N4909);
nor NOR4 (N5071, N5068, N241, N2266, N4374);
or OR2 (N5072, N5054, N3441);
nor NOR2 (N5073, N5065, N268);
and AND2 (N5074, N5063, N1075);
nand NAND2 (N5075, N5066, N1149);
xor XOR2 (N5076, N5074, N1271);
xor XOR2 (N5077, N5067, N577);
not NOT1 (N5078, N5044);
buf BUF1 (N5079, N5071);
buf BUF1 (N5080, N5072);
xor XOR2 (N5081, N5080, N531);
and AND2 (N5082, N5081, N5057);
not NOT1 (N5083, N5053);
or OR4 (N5084, N5082, N2376, N3661, N283);
xor XOR2 (N5085, N5076, N113);
nor NOR3 (N5086, N5083, N677, N2038);
buf BUF1 (N5087, N5085);
or OR4 (N5088, N5075, N1557, N735, N467);
nand NAND4 (N5089, N5079, N1629, N605, N2072);
or OR2 (N5090, N5070, N2086);
not NOT1 (N5091, N5069);
nor NOR3 (N5092, N5090, N3149, N3237);
and AND3 (N5093, N5084, N186, N3943);
and AND3 (N5094, N5073, N3356, N4673);
nand NAND2 (N5095, N5086, N4713);
not NOT1 (N5096, N5095);
nor NOR3 (N5097, N5094, N4276, N2736);
xor XOR2 (N5098, N5089, N1905);
not NOT1 (N5099, N5092);
xor XOR2 (N5100, N5096, N3898);
nand NAND4 (N5101, N5078, N4050, N2436, N2352);
or OR4 (N5102, N5088, N2041, N3983, N4898);
xor XOR2 (N5103, N5098, N4771);
not NOT1 (N5104, N5102);
not NOT1 (N5105, N5091);
not NOT1 (N5106, N5099);
buf BUF1 (N5107, N5101);
nor NOR3 (N5108, N5106, N3304, N694);
or OR4 (N5109, N5107, N4817, N440, N2006);
buf BUF1 (N5110, N5108);
or OR3 (N5111, N5087, N2910, N387);
and AND3 (N5112, N5104, N4908, N1319);
nor NOR2 (N5113, N5097, N2225);
nand NAND4 (N5114, N5100, N1636, N4286, N568);
buf BUF1 (N5115, N5114);
nand NAND2 (N5116, N5111, N3503);
or OR4 (N5117, N5115, N678, N2378, N3489);
nand NAND4 (N5118, N5112, N4634, N2061, N2495);
xor XOR2 (N5119, N5113, N2159);
and AND4 (N5120, N5110, N1812, N1650, N2688);
not NOT1 (N5121, N5119);
buf BUF1 (N5122, N5077);
xor XOR2 (N5123, N5122, N4036);
or OR3 (N5124, N5116, N545, N72);
or OR3 (N5125, N5123, N3845, N4755);
xor XOR2 (N5126, N5103, N1877);
nand NAND3 (N5127, N5121, N1281, N2456);
or OR2 (N5128, N5120, N2337);
or OR4 (N5129, N5117, N804, N3449, N1191);
xor XOR2 (N5130, N5109, N1708);
or OR3 (N5131, N5126, N1360, N847);
not NOT1 (N5132, N5131);
and AND4 (N5133, N5128, N3383, N4889, N1723);
nor NOR3 (N5134, N5130, N3629, N2116);
and AND3 (N5135, N5132, N3390, N2560);
and AND3 (N5136, N5134, N2946, N777);
xor XOR2 (N5137, N5136, N3550);
nand NAND2 (N5138, N5127, N227);
buf BUF1 (N5139, N5105);
or OR2 (N5140, N5133, N3628);
or OR3 (N5141, N5140, N2811, N1130);
buf BUF1 (N5142, N5137);
buf BUF1 (N5143, N5139);
and AND2 (N5144, N5143, N3085);
or OR4 (N5145, N5118, N2993, N1986, N2406);
xor XOR2 (N5146, N5125, N2605);
nor NOR3 (N5147, N5142, N4838, N921);
or OR2 (N5148, N5093, N1576);
or OR4 (N5149, N5138, N4363, N4755, N4957);
nand NAND4 (N5150, N5145, N4138, N2787, N957);
nor NOR3 (N5151, N5129, N3412, N4196);
or OR2 (N5152, N5147, N2108);
nor NOR3 (N5153, N5135, N830, N2469);
nor NOR4 (N5154, N5124, N1637, N3974, N2033);
not NOT1 (N5155, N5153);
or OR3 (N5156, N5150, N4188, N4353);
nor NOR2 (N5157, N5141, N2087);
nor NOR4 (N5158, N5146, N2366, N4426, N2221);
and AND2 (N5159, N5148, N4430);
buf BUF1 (N5160, N5156);
nor NOR4 (N5161, N5152, N4454, N2267, N3438);
not NOT1 (N5162, N5161);
nand NAND2 (N5163, N5155, N2212);
nand NAND2 (N5164, N5144, N1870);
buf BUF1 (N5165, N5160);
xor XOR2 (N5166, N5149, N1612);
not NOT1 (N5167, N5164);
nor NOR4 (N5168, N5154, N4474, N124, N22);
buf BUF1 (N5169, N5159);
xor XOR2 (N5170, N5157, N3812);
or OR4 (N5171, N5166, N1846, N640, N3577);
or OR2 (N5172, N5151, N3060);
xor XOR2 (N5173, N5165, N2921);
buf BUF1 (N5174, N5168);
buf BUF1 (N5175, N5173);
nor NOR2 (N5176, N5172, N2408);
nand NAND3 (N5177, N5169, N4491, N1382);
and AND4 (N5178, N5177, N221, N2536, N1263);
nor NOR2 (N5179, N5175, N2846);
xor XOR2 (N5180, N5162, N989);
or OR2 (N5181, N5167, N4632);
not NOT1 (N5182, N5158);
xor XOR2 (N5183, N5179, N4766);
or OR4 (N5184, N5178, N991, N1149, N2127);
nand NAND2 (N5185, N5174, N1000);
buf BUF1 (N5186, N5170);
xor XOR2 (N5187, N5181, N4733);
nand NAND4 (N5188, N5176, N5027, N1567, N2897);
and AND3 (N5189, N5184, N3919, N3732);
nand NAND2 (N5190, N5189, N5065);
buf BUF1 (N5191, N5171);
or OR4 (N5192, N5180, N3055, N4442, N1427);
buf BUF1 (N5193, N5191);
buf BUF1 (N5194, N5187);
and AND4 (N5195, N5185, N622, N1369, N3399);
not NOT1 (N5196, N5182);
or OR2 (N5197, N5186, N3935);
not NOT1 (N5198, N5183);
not NOT1 (N5199, N5195);
not NOT1 (N5200, N5163);
xor XOR2 (N5201, N5200, N984);
buf BUF1 (N5202, N5194);
and AND3 (N5203, N5196, N2475, N1087);
not NOT1 (N5204, N5203);
or OR3 (N5205, N5193, N2615, N558);
or OR3 (N5206, N5201, N4369, N1439);
buf BUF1 (N5207, N5192);
not NOT1 (N5208, N5198);
xor XOR2 (N5209, N5207, N2703);
xor XOR2 (N5210, N5208, N1271);
or OR4 (N5211, N5197, N568, N2607, N1625);
nor NOR2 (N5212, N5190, N2105);
or OR3 (N5213, N5211, N1338, N3781);
buf BUF1 (N5214, N5204);
nand NAND4 (N5215, N5213, N4568, N1647, N3530);
nor NOR4 (N5216, N5205, N3923, N2758, N4524);
nand NAND4 (N5217, N5202, N1795, N1160, N65);
or OR3 (N5218, N5216, N1916, N2169);
or OR2 (N5219, N5210, N3608);
not NOT1 (N5220, N5218);
nor NOR4 (N5221, N5209, N1950, N4765, N2682);
buf BUF1 (N5222, N5219);
or OR3 (N5223, N5188, N4324, N2898);
not NOT1 (N5224, N5199);
not NOT1 (N5225, N5221);
buf BUF1 (N5226, N5225);
xor XOR2 (N5227, N5226, N180);
or OR3 (N5228, N5215, N4821, N2524);
nand NAND4 (N5229, N5217, N1668, N4987, N5181);
and AND3 (N5230, N5229, N1533, N3168);
nand NAND2 (N5231, N5206, N2766);
not NOT1 (N5232, N5220);
not NOT1 (N5233, N5227);
or OR3 (N5234, N5224, N714, N4068);
and AND2 (N5235, N5212, N4269);
xor XOR2 (N5236, N5222, N1796);
nand NAND3 (N5237, N5231, N1293, N172);
buf BUF1 (N5238, N5223);
nor NOR4 (N5239, N5214, N2824, N895, N191);
or OR4 (N5240, N5228, N3854, N722, N1867);
buf BUF1 (N5241, N5234);
and AND4 (N5242, N5236, N1805, N7, N1541);
xor XOR2 (N5243, N5240, N4778);
or OR4 (N5244, N5237, N1754, N4178, N991);
not NOT1 (N5245, N5239);
and AND2 (N5246, N5241, N3629);
nand NAND4 (N5247, N5245, N4517, N3791, N1978);
or OR4 (N5248, N5238, N3860, N247, N3559);
buf BUF1 (N5249, N5248);
nand NAND3 (N5250, N5242, N3605, N4665);
and AND4 (N5251, N5232, N3084, N288, N1872);
nor NOR4 (N5252, N5235, N621, N1656, N2500);
buf BUF1 (N5253, N5246);
and AND4 (N5254, N5253, N3920, N1044, N2461);
not NOT1 (N5255, N5250);
and AND3 (N5256, N5233, N686, N4033);
or OR4 (N5257, N5243, N3708, N2200, N4057);
not NOT1 (N5258, N5257);
xor XOR2 (N5259, N5256, N313);
buf BUF1 (N5260, N5251);
or OR2 (N5261, N5259, N1305);
buf BUF1 (N5262, N5230);
xor XOR2 (N5263, N5249, N661);
buf BUF1 (N5264, N5263);
not NOT1 (N5265, N5255);
buf BUF1 (N5266, N5265);
nor NOR3 (N5267, N5258, N2934, N918);
or OR4 (N5268, N5244, N3384, N4769, N2659);
nand NAND3 (N5269, N5264, N3798, N22);
nand NAND3 (N5270, N5266, N1242, N2352);
nand NAND4 (N5271, N5252, N1358, N2452, N4020);
and AND4 (N5272, N5267, N2723, N389, N3779);
buf BUF1 (N5273, N5269);
nor NOR2 (N5274, N5261, N3621);
nor NOR4 (N5275, N5270, N1453, N3168, N1273);
or OR4 (N5276, N5247, N1918, N5249, N5121);
not NOT1 (N5277, N5276);
nor NOR3 (N5278, N5271, N1859, N763);
or OR3 (N5279, N5260, N1926, N2017);
nor NOR2 (N5280, N5262, N936);
buf BUF1 (N5281, N5254);
xor XOR2 (N5282, N5278, N1159);
buf BUF1 (N5283, N5275);
and AND3 (N5284, N5283, N5077, N1117);
nand NAND4 (N5285, N5268, N1364, N3692, N1136);
nand NAND4 (N5286, N5272, N1452, N2357, N5103);
nor NOR4 (N5287, N5282, N3647, N320, N2692);
xor XOR2 (N5288, N5285, N1771);
or OR4 (N5289, N5277, N2097, N4920, N1282);
nor NOR4 (N5290, N5289, N4904, N2412, N1814);
buf BUF1 (N5291, N5280);
not NOT1 (N5292, N5284);
nand NAND2 (N5293, N5291, N3920);
buf BUF1 (N5294, N5287);
not NOT1 (N5295, N5281);
nor NOR2 (N5296, N5288, N3765);
nand NAND3 (N5297, N5296, N4345, N3106);
not NOT1 (N5298, N5293);
not NOT1 (N5299, N5298);
not NOT1 (N5300, N5292);
and AND4 (N5301, N5279, N3224, N3325, N783);
nand NAND3 (N5302, N5273, N1728, N1486);
and AND2 (N5303, N5274, N4183);
nand NAND3 (N5304, N5300, N2458, N3387);
buf BUF1 (N5305, N5299);
buf BUF1 (N5306, N5295);
nor NOR3 (N5307, N5306, N1898, N4628);
xor XOR2 (N5308, N5301, N5073);
not NOT1 (N5309, N5308);
xor XOR2 (N5310, N5302, N2652);
buf BUF1 (N5311, N5310);
nor NOR4 (N5312, N5305, N3008, N1199, N1483);
not NOT1 (N5313, N5312);
not NOT1 (N5314, N5309);
buf BUF1 (N5315, N5311);
not NOT1 (N5316, N5314);
or OR4 (N5317, N5307, N1111, N5005, N2496);
not NOT1 (N5318, N5303);
nand NAND4 (N5319, N5290, N4469, N4531, N4951);
and AND4 (N5320, N5304, N1358, N754, N3858);
nor NOR3 (N5321, N5320, N2023, N345);
not NOT1 (N5322, N5321);
not NOT1 (N5323, N5316);
not NOT1 (N5324, N5286);
not NOT1 (N5325, N5317);
nand NAND3 (N5326, N5297, N1100, N3289);
or OR4 (N5327, N5318, N4545, N774, N2999);
and AND3 (N5328, N5322, N1151, N2699);
nor NOR3 (N5329, N5294, N3724, N1728);
xor XOR2 (N5330, N5327, N5311);
buf BUF1 (N5331, N5313);
nor NOR3 (N5332, N5328, N5061, N2542);
or OR4 (N5333, N5325, N2044, N748, N2680);
xor XOR2 (N5334, N5330, N795);
buf BUF1 (N5335, N5331);
or OR2 (N5336, N5319, N4224);
or OR2 (N5337, N5323, N14);
nand NAND3 (N5338, N5335, N1810, N3604);
nor NOR3 (N5339, N5334, N4257, N3517);
not NOT1 (N5340, N5315);
xor XOR2 (N5341, N5339, N5005);
nor NOR4 (N5342, N5326, N5127, N482, N2216);
not NOT1 (N5343, N5338);
and AND3 (N5344, N5336, N3730, N1418);
xor XOR2 (N5345, N5324, N3738);
not NOT1 (N5346, N5332);
buf BUF1 (N5347, N5337);
nor NOR2 (N5348, N5329, N3348);
buf BUF1 (N5349, N5344);
nor NOR2 (N5350, N5341, N149);
buf BUF1 (N5351, N5346);
or OR3 (N5352, N5343, N1116, N3076);
not NOT1 (N5353, N5347);
and AND3 (N5354, N5352, N5295, N233);
buf BUF1 (N5355, N5333);
buf BUF1 (N5356, N5342);
and AND3 (N5357, N5353, N2064, N2164);
buf BUF1 (N5358, N5356);
and AND4 (N5359, N5340, N4517, N1233, N4264);
buf BUF1 (N5360, N5357);
nor NOR2 (N5361, N5349, N4456);
buf BUF1 (N5362, N5351);
xor XOR2 (N5363, N5348, N356);
not NOT1 (N5364, N5363);
nand NAND3 (N5365, N5345, N5060, N3364);
buf BUF1 (N5366, N5364);
and AND4 (N5367, N5350, N1939, N2817, N4635);
and AND4 (N5368, N5361, N2464, N2044, N3482);
and AND3 (N5369, N5359, N2306, N4364);
nand NAND3 (N5370, N5360, N2340, N3745);
not NOT1 (N5371, N5358);
nor NOR3 (N5372, N5355, N3752, N970);
nor NOR3 (N5373, N5372, N850, N2753);
nand NAND2 (N5374, N5369, N4490);
and AND3 (N5375, N5365, N3016, N3112);
or OR4 (N5376, N5374, N421, N3018, N2979);
nor NOR4 (N5377, N5367, N4744, N4185, N3096);
nor NOR4 (N5378, N5377, N1427, N141, N3652);
and AND2 (N5379, N5373, N2027);
nor NOR2 (N5380, N5368, N4522);
nor NOR3 (N5381, N5380, N2301, N4050);
buf BUF1 (N5382, N5381);
and AND2 (N5383, N5362, N664);
or OR4 (N5384, N5376, N3797, N2207, N4519);
nor NOR4 (N5385, N5379, N436, N4702, N3237);
not NOT1 (N5386, N5371);
and AND2 (N5387, N5375, N2262);
or OR4 (N5388, N5354, N3941, N896, N1908);
or OR4 (N5389, N5385, N5094, N4694, N1124);
not NOT1 (N5390, N5389);
nor NOR3 (N5391, N5388, N1563, N4543);
buf BUF1 (N5392, N5384);
nand NAND2 (N5393, N5370, N1219);
nor NOR4 (N5394, N5382, N4832, N675, N188);
or OR3 (N5395, N5392, N1263, N4524);
xor XOR2 (N5396, N5378, N2779);
or OR4 (N5397, N5386, N3154, N3311, N3569);
xor XOR2 (N5398, N5393, N1846);
or OR3 (N5399, N5391, N402, N2155);
and AND3 (N5400, N5366, N202, N613);
nand NAND3 (N5401, N5400, N1108, N4380);
not NOT1 (N5402, N5383);
and AND4 (N5403, N5399, N1354, N3453, N5166);
buf BUF1 (N5404, N5403);
not NOT1 (N5405, N5398);
or OR3 (N5406, N5404, N366, N906);
or OR2 (N5407, N5406, N1778);
nand NAND4 (N5408, N5390, N738, N2578, N3041);
xor XOR2 (N5409, N5397, N2468);
or OR2 (N5410, N5394, N2866);
not NOT1 (N5411, N5409);
or OR4 (N5412, N5408, N344, N4343, N2559);
nand NAND2 (N5413, N5396, N2108);
nor NOR3 (N5414, N5412, N5375, N124);
nand NAND4 (N5415, N5413, N105, N1465, N283);
and AND2 (N5416, N5402, N2463);
xor XOR2 (N5417, N5387, N2455);
buf BUF1 (N5418, N5401);
buf BUF1 (N5419, N5395);
not NOT1 (N5420, N5411);
not NOT1 (N5421, N5415);
or OR2 (N5422, N5421, N386);
not NOT1 (N5423, N5419);
not NOT1 (N5424, N5405);
nand NAND3 (N5425, N5416, N2918, N1356);
and AND2 (N5426, N5424, N752);
buf BUF1 (N5427, N5423);
not NOT1 (N5428, N5417);
and AND3 (N5429, N5427, N3512, N1654);
not NOT1 (N5430, N5422);
xor XOR2 (N5431, N5429, N2568);
nor NOR3 (N5432, N5430, N2476, N3272);
xor XOR2 (N5433, N5432, N431);
nand NAND3 (N5434, N5410, N1257, N672);
nand NAND2 (N5435, N5425, N5075);
buf BUF1 (N5436, N5431);
nand NAND4 (N5437, N5426, N1379, N2450, N758);
buf BUF1 (N5438, N5407);
xor XOR2 (N5439, N5436, N4613);
buf BUF1 (N5440, N5437);
nor NOR4 (N5441, N5420, N782, N2847, N5331);
and AND3 (N5442, N5433, N3736, N4845);
nor NOR3 (N5443, N5442, N3247, N2434);
xor XOR2 (N5444, N5439, N4500);
nor NOR4 (N5445, N5434, N1802, N37, N2341);
nor NOR2 (N5446, N5444, N1228);
buf BUF1 (N5447, N5435);
or OR2 (N5448, N5418, N1369);
xor XOR2 (N5449, N5445, N1516);
or OR2 (N5450, N5449, N204);
or OR4 (N5451, N5428, N4958, N824, N3679);
buf BUF1 (N5452, N5443);
and AND3 (N5453, N5414, N4415, N1990);
buf BUF1 (N5454, N5446);
and AND3 (N5455, N5438, N1521, N286);
or OR4 (N5456, N5455, N3931, N2535, N1618);
or OR2 (N5457, N5447, N5206);
nand NAND3 (N5458, N5451, N2248, N4949);
xor XOR2 (N5459, N5441, N4671);
buf BUF1 (N5460, N5450);
not NOT1 (N5461, N5453);
nand NAND3 (N5462, N5440, N231, N62);
xor XOR2 (N5463, N5454, N4804);
not NOT1 (N5464, N5457);
xor XOR2 (N5465, N5463, N2647);
or OR2 (N5466, N5460, N1008);
nor NOR4 (N5467, N5466, N3891, N65, N3218);
nand NAND2 (N5468, N5448, N3859);
nor NOR3 (N5469, N5458, N4062, N4596);
nor NOR3 (N5470, N5452, N3767, N2075);
nor NOR3 (N5471, N5459, N4407, N1270);
not NOT1 (N5472, N5471);
nor NOR4 (N5473, N5461, N2408, N2882, N38);
buf BUF1 (N5474, N5473);
or OR3 (N5475, N5474, N3875, N2133);
and AND4 (N5476, N5475, N328, N4961, N4974);
xor XOR2 (N5477, N5464, N1939);
buf BUF1 (N5478, N5467);
nand NAND4 (N5479, N5456, N1125, N2554, N4077);
xor XOR2 (N5480, N5469, N967);
not NOT1 (N5481, N5479);
nor NOR2 (N5482, N5465, N2113);
buf BUF1 (N5483, N5481);
not NOT1 (N5484, N5483);
not NOT1 (N5485, N5478);
nand NAND4 (N5486, N5476, N1469, N1131, N4371);
xor XOR2 (N5487, N5477, N3093);
or OR2 (N5488, N5482, N159);
nand NAND4 (N5489, N5487, N3403, N3401, N5376);
nand NAND4 (N5490, N5468, N2570, N2140, N262);
or OR4 (N5491, N5488, N4991, N187, N370);
nor NOR2 (N5492, N5484, N2142);
and AND2 (N5493, N5480, N5458);
buf BUF1 (N5494, N5492);
nor NOR3 (N5495, N5489, N1735, N2439);
and AND2 (N5496, N5462, N1090);
buf BUF1 (N5497, N5472);
and AND2 (N5498, N5486, N3640);
nor NOR2 (N5499, N5496, N1542);
not NOT1 (N5500, N5498);
nand NAND2 (N5501, N5497, N624);
buf BUF1 (N5502, N5494);
xor XOR2 (N5503, N5490, N3332);
and AND2 (N5504, N5491, N3427);
not NOT1 (N5505, N5503);
nand NAND4 (N5506, N5499, N4700, N3239, N2129);
nand NAND3 (N5507, N5485, N5161, N4382);
and AND3 (N5508, N5505, N3636, N4504);
nand NAND2 (N5509, N5500, N1229);
and AND3 (N5510, N5504, N3739, N3699);
buf BUF1 (N5511, N5495);
buf BUF1 (N5512, N5493);
and AND2 (N5513, N5470, N1239);
not NOT1 (N5514, N5512);
and AND3 (N5515, N5509, N1383, N4120);
nand NAND3 (N5516, N5506, N423, N3689);
nor NOR4 (N5517, N5508, N1101, N442, N800);
not NOT1 (N5518, N5502);
and AND2 (N5519, N5514, N566);
nor NOR4 (N5520, N5517, N5193, N649, N5222);
xor XOR2 (N5521, N5511, N1164);
or OR3 (N5522, N5520, N1719, N3189);
not NOT1 (N5523, N5516);
nand NAND2 (N5524, N5521, N2726);
nor NOR3 (N5525, N5518, N2881, N1255);
not NOT1 (N5526, N5510);
or OR2 (N5527, N5513, N1858);
not NOT1 (N5528, N5523);
and AND4 (N5529, N5522, N4291, N2763, N3913);
nor NOR2 (N5530, N5515, N4449);
or OR4 (N5531, N5529, N5402, N3024, N1150);
nand NAND2 (N5532, N5519, N1427);
nand NAND2 (N5533, N5501, N2946);
nor NOR3 (N5534, N5526, N1676, N2932);
nor NOR4 (N5535, N5532, N290, N2848, N5429);
buf BUF1 (N5536, N5528);
or OR3 (N5537, N5531, N1655, N3841);
or OR2 (N5538, N5524, N1149);
or OR3 (N5539, N5535, N2131, N4313);
and AND2 (N5540, N5539, N1897);
not NOT1 (N5541, N5530);
xor XOR2 (N5542, N5525, N2660);
xor XOR2 (N5543, N5538, N3150);
xor XOR2 (N5544, N5537, N4946);
and AND4 (N5545, N5540, N5426, N955, N3502);
xor XOR2 (N5546, N5542, N3963);
nand NAND2 (N5547, N5507, N3276);
buf BUF1 (N5548, N5547);
nand NAND4 (N5549, N5545, N94, N91, N846);
xor XOR2 (N5550, N5546, N3024);
buf BUF1 (N5551, N5533);
nand NAND2 (N5552, N5550, N2106);
nand NAND3 (N5553, N5548, N2642, N2670);
xor XOR2 (N5554, N5543, N5186);
not NOT1 (N5555, N5553);
buf BUF1 (N5556, N5554);
nand NAND2 (N5557, N5527, N1011);
nor NOR3 (N5558, N5536, N2665, N3215);
nor NOR3 (N5559, N5557, N5511, N2833);
nor NOR3 (N5560, N5555, N1298, N4124);
or OR2 (N5561, N5552, N1609);
buf BUF1 (N5562, N5541);
nor NOR2 (N5563, N5559, N603);
buf BUF1 (N5564, N5558);
and AND2 (N5565, N5534, N3455);
buf BUF1 (N5566, N5564);
not NOT1 (N5567, N5562);
and AND2 (N5568, N5561, N1400);
nor NOR2 (N5569, N5566, N968);
and AND4 (N5570, N5565, N666, N1578, N3952);
or OR2 (N5571, N5568, N1865);
buf BUF1 (N5572, N5571);
and AND4 (N5573, N5551, N1510, N675, N179);
or OR2 (N5574, N5560, N1228);
xor XOR2 (N5575, N5563, N4760);
and AND2 (N5576, N5572, N5119);
and AND2 (N5577, N5576, N242);
or OR2 (N5578, N5577, N5354);
not NOT1 (N5579, N5544);
and AND2 (N5580, N5556, N1393);
nand NAND3 (N5581, N5580, N2435, N277);
xor XOR2 (N5582, N5574, N428);
and AND4 (N5583, N5575, N3367, N3169, N4460);
not NOT1 (N5584, N5569);
xor XOR2 (N5585, N5573, N3736);
or OR3 (N5586, N5582, N1134, N1813);
not NOT1 (N5587, N5570);
or OR2 (N5588, N5587, N3095);
nor NOR4 (N5589, N5578, N4146, N4046, N1792);
xor XOR2 (N5590, N5581, N3052);
buf BUF1 (N5591, N5567);
not NOT1 (N5592, N5584);
buf BUF1 (N5593, N5549);
xor XOR2 (N5594, N5593, N5196);
not NOT1 (N5595, N5592);
nand NAND4 (N5596, N5594, N529, N1608, N3814);
and AND3 (N5597, N5588, N4065, N124);
nand NAND3 (N5598, N5597, N4788, N835);
or OR2 (N5599, N5595, N4423);
nor NOR2 (N5600, N5599, N3319);
and AND4 (N5601, N5590, N1566, N2334, N4091);
not NOT1 (N5602, N5583);
nand NAND4 (N5603, N5591, N3359, N2220, N3899);
nand NAND3 (N5604, N5585, N1928, N3591);
buf BUF1 (N5605, N5600);
nor NOR4 (N5606, N5589, N1806, N1934, N2605);
xor XOR2 (N5607, N5598, N2686);
xor XOR2 (N5608, N5603, N1628);
nand NAND3 (N5609, N5608, N3894, N5413);
and AND3 (N5610, N5605, N2384, N837);
buf BUF1 (N5611, N5602);
or OR2 (N5612, N5586, N3099);
and AND4 (N5613, N5579, N4132, N373, N49);
nor NOR3 (N5614, N5607, N2063, N5603);
not NOT1 (N5615, N5604);
or OR3 (N5616, N5606, N311, N990);
not NOT1 (N5617, N5613);
nor NOR4 (N5618, N5617, N667, N1871, N3491);
and AND4 (N5619, N5610, N3402, N1392, N1657);
xor XOR2 (N5620, N5601, N5280);
nor NOR2 (N5621, N5609, N1982);
buf BUF1 (N5622, N5618);
not NOT1 (N5623, N5619);
buf BUF1 (N5624, N5611);
nand NAND3 (N5625, N5614, N3785, N471);
nor NOR2 (N5626, N5622, N66);
nor NOR4 (N5627, N5620, N134, N628, N292);
and AND4 (N5628, N5621, N1721, N2390, N4873);
buf BUF1 (N5629, N5596);
nor NOR3 (N5630, N5625, N3218, N4567);
xor XOR2 (N5631, N5624, N1666);
xor XOR2 (N5632, N5612, N2176);
xor XOR2 (N5633, N5615, N5266);
buf BUF1 (N5634, N5631);
nor NOR3 (N5635, N5629, N5372, N5389);
xor XOR2 (N5636, N5633, N4159);
nand NAND3 (N5637, N5616, N5411, N4546);
and AND4 (N5638, N5636, N162, N1116, N1647);
xor XOR2 (N5639, N5626, N2288);
and AND2 (N5640, N5632, N2603);
nand NAND3 (N5641, N5634, N2503, N222);
nand NAND4 (N5642, N5638, N2867, N2553, N772);
buf BUF1 (N5643, N5639);
nor NOR3 (N5644, N5641, N2093, N2127);
nand NAND4 (N5645, N5642, N4020, N2516, N4159);
xor XOR2 (N5646, N5630, N5547);
nor NOR3 (N5647, N5643, N4934, N4964);
buf BUF1 (N5648, N5646);
or OR2 (N5649, N5628, N2402);
xor XOR2 (N5650, N5645, N3949);
not NOT1 (N5651, N5627);
nand NAND2 (N5652, N5651, N362);
nand NAND4 (N5653, N5647, N1915, N2200, N3657);
and AND2 (N5654, N5649, N1044);
or OR2 (N5655, N5650, N161);
nor NOR2 (N5656, N5655, N1895);
not NOT1 (N5657, N5648);
and AND3 (N5658, N5640, N5538, N5382);
nand NAND4 (N5659, N5623, N4203, N4060, N697);
nor NOR2 (N5660, N5653, N440);
nor NOR3 (N5661, N5660, N5419, N3177);
not NOT1 (N5662, N5635);
buf BUF1 (N5663, N5659);
buf BUF1 (N5664, N5661);
nand NAND4 (N5665, N5664, N343, N1865, N2213);
nor NOR4 (N5666, N5663, N861, N1064, N3968);
xor XOR2 (N5667, N5666, N924);
nor NOR4 (N5668, N5644, N3109, N4404, N941);
nand NAND3 (N5669, N5652, N405, N469);
or OR3 (N5670, N5637, N1039, N3657);
and AND4 (N5671, N5670, N3347, N4821, N2418);
or OR2 (N5672, N5667, N705);
nor NOR2 (N5673, N5656, N278);
not NOT1 (N5674, N5672);
buf BUF1 (N5675, N5674);
nor NOR4 (N5676, N5657, N3332, N4889, N861);
nor NOR4 (N5677, N5669, N3077, N2501, N92);
and AND4 (N5678, N5662, N1772, N1377, N1861);
nand NAND3 (N5679, N5654, N107, N1031);
nor NOR4 (N5680, N5677, N2187, N4419, N1955);
nand NAND2 (N5681, N5673, N2291);
or OR4 (N5682, N5680, N5429, N805, N4576);
xor XOR2 (N5683, N5658, N2664);
buf BUF1 (N5684, N5675);
or OR4 (N5685, N5682, N3555, N220, N745);
nand NAND4 (N5686, N5685, N2339, N246, N475);
xor XOR2 (N5687, N5681, N710);
and AND3 (N5688, N5665, N1872, N2262);
xor XOR2 (N5689, N5668, N2079);
and AND2 (N5690, N5684, N557);
nor NOR2 (N5691, N5686, N2699);
nor NOR4 (N5692, N5689, N4930, N5606, N3247);
not NOT1 (N5693, N5692);
xor XOR2 (N5694, N5690, N1764);
and AND3 (N5695, N5688, N861, N2996);
nor NOR4 (N5696, N5671, N3579, N5202, N429);
buf BUF1 (N5697, N5696);
not NOT1 (N5698, N5676);
buf BUF1 (N5699, N5693);
xor XOR2 (N5700, N5687, N2515);
and AND2 (N5701, N5679, N2148);
and AND3 (N5702, N5700, N745, N73);
or OR3 (N5703, N5694, N968, N2342);
nand NAND2 (N5704, N5691, N351);
buf BUF1 (N5705, N5699);
not NOT1 (N5706, N5678);
or OR2 (N5707, N5705, N809);
buf BUF1 (N5708, N5683);
xor XOR2 (N5709, N5698, N978);
nor NOR3 (N5710, N5704, N5343, N5092);
nand NAND4 (N5711, N5701, N1761, N1204, N1085);
buf BUF1 (N5712, N5708);
or OR2 (N5713, N5702, N5053);
not NOT1 (N5714, N5712);
nand NAND2 (N5715, N5713, N821);
not NOT1 (N5716, N5707);
nand NAND4 (N5717, N5703, N612, N3810, N1307);
xor XOR2 (N5718, N5695, N1990);
and AND3 (N5719, N5715, N1348, N2763);
xor XOR2 (N5720, N5717, N3278);
buf BUF1 (N5721, N5718);
and AND3 (N5722, N5697, N3659, N503);
xor XOR2 (N5723, N5719, N1114);
nand NAND4 (N5724, N5723, N825, N1873, N768);
buf BUF1 (N5725, N5714);
and AND3 (N5726, N5709, N4004, N1779);
not NOT1 (N5727, N5722);
not NOT1 (N5728, N5716);
nand NAND4 (N5729, N5720, N2612, N2370, N2623);
nand NAND4 (N5730, N5727, N1277, N4049, N4427);
buf BUF1 (N5731, N5710);
nor NOR3 (N5732, N5728, N4799, N3672);
nand NAND3 (N5733, N5726, N3091, N3981);
buf BUF1 (N5734, N5724);
buf BUF1 (N5735, N5731);
xor XOR2 (N5736, N5721, N4331);
buf BUF1 (N5737, N5730);
nand NAND2 (N5738, N5732, N4636);
nor NOR4 (N5739, N5734, N4992, N5719, N3479);
nor NOR2 (N5740, N5725, N982);
and AND3 (N5741, N5739, N298, N3127);
nor NOR4 (N5742, N5737, N4895, N4372, N1577);
and AND2 (N5743, N5735, N661);
xor XOR2 (N5744, N5706, N236);
xor XOR2 (N5745, N5711, N4609);
nand NAND4 (N5746, N5740, N1553, N1122, N2718);
xor XOR2 (N5747, N5746, N7);
nor NOR3 (N5748, N5736, N1814, N503);
nor NOR2 (N5749, N5742, N2533);
xor XOR2 (N5750, N5738, N2420);
xor XOR2 (N5751, N5741, N2593);
and AND3 (N5752, N5744, N1442, N802);
not NOT1 (N5753, N5748);
buf BUF1 (N5754, N5753);
not NOT1 (N5755, N5733);
xor XOR2 (N5756, N5750, N2219);
and AND3 (N5757, N5752, N4425, N4780);
nor NOR2 (N5758, N5756, N2902);
or OR3 (N5759, N5729, N1975, N213);
xor XOR2 (N5760, N5758, N4431);
or OR4 (N5761, N5757, N414, N893, N3588);
nor NOR4 (N5762, N5761, N4489, N2057, N1811);
or OR4 (N5763, N5745, N5003, N557, N5136);
not NOT1 (N5764, N5747);
or OR3 (N5765, N5759, N559, N3448);
not NOT1 (N5766, N5755);
or OR4 (N5767, N5764, N1279, N3037, N905);
or OR3 (N5768, N5765, N640, N3160);
xor XOR2 (N5769, N5768, N863);
buf BUF1 (N5770, N5749);
nand NAND4 (N5771, N5766, N2063, N3908, N757);
xor XOR2 (N5772, N5743, N249);
nor NOR3 (N5773, N5767, N1036, N779);
nor NOR4 (N5774, N5769, N3186, N4805, N472);
and AND3 (N5775, N5762, N3995, N1530);
or OR3 (N5776, N5773, N4504, N538);
nand NAND3 (N5777, N5771, N2633, N678);
or OR3 (N5778, N5754, N4083, N4137);
nand NAND2 (N5779, N5751, N5425);
buf BUF1 (N5780, N5775);
xor XOR2 (N5781, N5780, N2546);
or OR2 (N5782, N5778, N5533);
or OR2 (N5783, N5779, N259);
not NOT1 (N5784, N5777);
buf BUF1 (N5785, N5772);
nor NOR3 (N5786, N5760, N5673, N2264);
buf BUF1 (N5787, N5774);
not NOT1 (N5788, N5786);
nand NAND3 (N5789, N5776, N3029, N4490);
nand NAND3 (N5790, N5782, N2325, N3899);
nor NOR3 (N5791, N5787, N4382, N1486);
nor NOR3 (N5792, N5791, N319, N4541);
nor NOR4 (N5793, N5792, N2513, N4304, N4341);
xor XOR2 (N5794, N5789, N5293);
nand NAND4 (N5795, N5790, N2506, N3578, N4319);
not NOT1 (N5796, N5795);
nand NAND3 (N5797, N5770, N5700, N2767);
nor NOR4 (N5798, N5785, N3108, N1894, N1375);
nand NAND3 (N5799, N5797, N2409, N4271);
and AND3 (N5800, N5788, N5065, N3589);
nand NAND4 (N5801, N5783, N1946, N3705, N1974);
and AND2 (N5802, N5800, N1366);
buf BUF1 (N5803, N5801);
buf BUF1 (N5804, N5796);
xor XOR2 (N5805, N5802, N1519);
or OR4 (N5806, N5763, N2224, N1556, N3810);
buf BUF1 (N5807, N5803);
buf BUF1 (N5808, N5805);
buf BUF1 (N5809, N5793);
not NOT1 (N5810, N5807);
nor NOR2 (N5811, N5781, N2966);
nor NOR2 (N5812, N5809, N1719);
or OR3 (N5813, N5784, N2637, N3171);
buf BUF1 (N5814, N5794);
not NOT1 (N5815, N5804);
not NOT1 (N5816, N5798);
or OR3 (N5817, N5806, N1916, N694);
nand NAND3 (N5818, N5812, N2985, N694);
or OR2 (N5819, N5808, N3820);
and AND4 (N5820, N5816, N1945, N2568, N5445);
or OR2 (N5821, N5810, N5484);
xor XOR2 (N5822, N5811, N656);
and AND2 (N5823, N5820, N5637);
or OR2 (N5824, N5817, N1443);
not NOT1 (N5825, N5799);
nand NAND2 (N5826, N5813, N5415);
nand NAND2 (N5827, N5823, N2703);
not NOT1 (N5828, N5824);
not NOT1 (N5829, N5815);
xor XOR2 (N5830, N5827, N3097);
or OR3 (N5831, N5825, N2047, N2452);
nor NOR2 (N5832, N5829, N3688);
and AND4 (N5833, N5821, N2949, N4302, N1464);
nand NAND4 (N5834, N5833, N4335, N5474, N4926);
not NOT1 (N5835, N5830);
or OR2 (N5836, N5834, N5049);
buf BUF1 (N5837, N5832);
and AND4 (N5838, N5831, N72, N4643, N1073);
xor XOR2 (N5839, N5826, N3833);
buf BUF1 (N5840, N5836);
nand NAND4 (N5841, N5839, N2857, N3978, N1302);
not NOT1 (N5842, N5814);
nor NOR4 (N5843, N5837, N2831, N716, N3584);
or OR2 (N5844, N5840, N1341);
or OR2 (N5845, N5818, N3309);
or OR3 (N5846, N5843, N971, N5760);
nor NOR4 (N5847, N5838, N3145, N892, N2428);
not NOT1 (N5848, N5828);
not NOT1 (N5849, N5844);
xor XOR2 (N5850, N5849, N2665);
nand NAND4 (N5851, N5846, N446, N4069, N2774);
and AND2 (N5852, N5842, N3415);
not NOT1 (N5853, N5852);
nand NAND3 (N5854, N5850, N3792, N1588);
buf BUF1 (N5855, N5819);
and AND3 (N5856, N5855, N688, N5076);
or OR4 (N5857, N5822, N5115, N239, N2268);
and AND4 (N5858, N5847, N5190, N3514, N1344);
xor XOR2 (N5859, N5835, N3360);
nand NAND4 (N5860, N5851, N5554, N1167, N5334);
not NOT1 (N5861, N5841);
nand NAND4 (N5862, N5845, N3306, N2558, N732);
and AND2 (N5863, N5859, N2282);
and AND4 (N5864, N5857, N1975, N2446, N5415);
or OR2 (N5865, N5854, N2720);
not NOT1 (N5866, N5858);
nor NOR4 (N5867, N5861, N4421, N2163, N5550);
and AND3 (N5868, N5867, N2886, N5436);
and AND3 (N5869, N5864, N2253, N3794);
or OR2 (N5870, N5853, N4626);
nor NOR2 (N5871, N5856, N191);
nor NOR2 (N5872, N5865, N5808);
buf BUF1 (N5873, N5871);
and AND3 (N5874, N5862, N921, N5729);
and AND3 (N5875, N5873, N2139, N616);
nor NOR2 (N5876, N5866, N5225);
xor XOR2 (N5877, N5875, N2800);
nor NOR4 (N5878, N5872, N3645, N797, N917);
nor NOR4 (N5879, N5878, N209, N5303, N982);
not NOT1 (N5880, N5877);
buf BUF1 (N5881, N5874);
nand NAND3 (N5882, N5881, N2417, N1829);
and AND4 (N5883, N5882, N5485, N1367, N4867);
nor NOR4 (N5884, N5860, N5815, N626, N4451);
nor NOR3 (N5885, N5883, N2868, N1937);
not NOT1 (N5886, N5848);
buf BUF1 (N5887, N5879);
or OR4 (N5888, N5869, N4063, N4561, N2752);
or OR2 (N5889, N5868, N4748);
nor NOR2 (N5890, N5880, N2149);
or OR2 (N5891, N5876, N3780);
not NOT1 (N5892, N5890);
nor NOR2 (N5893, N5891, N5651);
nand NAND4 (N5894, N5870, N481, N5668, N3164);
buf BUF1 (N5895, N5888);
xor XOR2 (N5896, N5863, N2537);
nand NAND3 (N5897, N5889, N4006, N1948);
or OR2 (N5898, N5895, N3931);
xor XOR2 (N5899, N5896, N3954);
xor XOR2 (N5900, N5898, N652);
nor NOR2 (N5901, N5885, N1363);
nand NAND2 (N5902, N5897, N2640);
nand NAND2 (N5903, N5887, N4314);
not NOT1 (N5904, N5903);
and AND2 (N5905, N5901, N916);
buf BUF1 (N5906, N5894);
and AND3 (N5907, N5893, N5671, N2141);
nand NAND3 (N5908, N5907, N166, N3669);
not NOT1 (N5909, N5886);
buf BUF1 (N5910, N5908);
nor NOR4 (N5911, N5900, N909, N1820, N4919);
not NOT1 (N5912, N5902);
and AND4 (N5913, N5904, N831, N5781, N2504);
nand NAND2 (N5914, N5892, N5098);
xor XOR2 (N5915, N5905, N2836);
or OR2 (N5916, N5911, N4214);
buf BUF1 (N5917, N5899);
nor NOR3 (N5918, N5884, N1490, N3227);
nor NOR3 (N5919, N5915, N1754, N2587);
and AND3 (N5920, N5913, N162, N12);
nor NOR2 (N5921, N5914, N5405);
nor NOR3 (N5922, N5920, N2291, N2908);
and AND3 (N5923, N5912, N3274, N3355);
xor XOR2 (N5924, N5919, N3811);
buf BUF1 (N5925, N5923);
buf BUF1 (N5926, N5922);
buf BUF1 (N5927, N5921);
buf BUF1 (N5928, N5918);
nor NOR3 (N5929, N5927, N2902, N291);
not NOT1 (N5930, N5924);
xor XOR2 (N5931, N5929, N3849);
buf BUF1 (N5932, N5917);
nor NOR3 (N5933, N5930, N636, N1299);
buf BUF1 (N5934, N5931);
nor NOR2 (N5935, N5928, N2162);
nand NAND4 (N5936, N5916, N1220, N204, N5933);
or OR2 (N5937, N889, N3180);
nand NAND4 (N5938, N5934, N91, N5307, N689);
or OR2 (N5939, N5926, N2367);
or OR3 (N5940, N5939, N4374, N5615);
nor NOR3 (N5941, N5910, N1018, N3005);
nand NAND2 (N5942, N5938, N1020);
and AND4 (N5943, N5942, N1035, N122, N645);
buf BUF1 (N5944, N5940);
and AND4 (N5945, N5943, N2891, N2213, N1620);
nor NOR3 (N5946, N5944, N4348, N502);
buf BUF1 (N5947, N5945);
or OR2 (N5948, N5906, N773);
buf BUF1 (N5949, N5909);
xor XOR2 (N5950, N5949, N1949);
nor NOR4 (N5951, N5947, N4024, N3057, N1092);
and AND3 (N5952, N5946, N1622, N475);
xor XOR2 (N5953, N5925, N5768);
buf BUF1 (N5954, N5952);
and AND2 (N5955, N5936, N4465);
not NOT1 (N5956, N5953);
xor XOR2 (N5957, N5956, N2366);
or OR3 (N5958, N5950, N2035, N931);
and AND4 (N5959, N5948, N2362, N2184, N3265);
xor XOR2 (N5960, N5954, N674);
or OR3 (N5961, N5957, N4736, N1199);
or OR3 (N5962, N5951, N2436, N5033);
or OR2 (N5963, N5962, N2322);
or OR3 (N5964, N5935, N711, N2502);
xor XOR2 (N5965, N5932, N2951);
nor NOR2 (N5966, N5937, N1475);
nor NOR3 (N5967, N5964, N1206, N1353);
or OR2 (N5968, N5960, N3449);
and AND3 (N5969, N5955, N5289, N345);
buf BUF1 (N5970, N5965);
buf BUF1 (N5971, N5968);
buf BUF1 (N5972, N5970);
and AND2 (N5973, N5967, N923);
or OR4 (N5974, N5973, N2545, N2674, N3553);
and AND4 (N5975, N5958, N1297, N5484, N2192);
nor NOR2 (N5976, N5974, N282);
and AND2 (N5977, N5966, N4879);
nand NAND3 (N5978, N5959, N319, N3332);
nor NOR2 (N5979, N5978, N1826);
and AND2 (N5980, N5963, N3583);
nor NOR2 (N5981, N5979, N1756);
and AND2 (N5982, N5971, N969);
not NOT1 (N5983, N5981);
or OR3 (N5984, N5972, N261, N2050);
xor XOR2 (N5985, N5983, N2153);
and AND2 (N5986, N5982, N164);
or OR4 (N5987, N5976, N2364, N5524, N471);
nor NOR3 (N5988, N5985, N4521, N1826);
nor NOR2 (N5989, N5941, N1571);
not NOT1 (N5990, N5988);
nand NAND2 (N5991, N5987, N1306);
xor XOR2 (N5992, N5975, N4400);
xor XOR2 (N5993, N5986, N455);
nor NOR3 (N5994, N5977, N1843, N4062);
buf BUF1 (N5995, N5980);
not NOT1 (N5996, N5990);
nand NAND2 (N5997, N5992, N355);
xor XOR2 (N5998, N5969, N3255);
nand NAND4 (N5999, N5961, N3469, N3887, N4173);
xor XOR2 (N6000, N5993, N4042);
xor XOR2 (N6001, N5997, N4615);
nand NAND3 (N6002, N5994, N4815, N4534);
and AND4 (N6003, N6000, N1987, N3408, N3661);
not NOT1 (N6004, N5989);
nand NAND3 (N6005, N6002, N3141, N2027);
or OR3 (N6006, N6005, N1205, N5027);
nor NOR4 (N6007, N6004, N1753, N4130, N437);
not NOT1 (N6008, N5984);
not NOT1 (N6009, N6003);
nor NOR4 (N6010, N5996, N840, N4745, N4373);
nand NAND2 (N6011, N6009, N4177);
and AND3 (N6012, N6001, N1679, N2055);
or OR3 (N6013, N6010, N3917, N4628);
and AND2 (N6014, N6007, N1996);
or OR4 (N6015, N5995, N4532, N3778, N2823);
nand NAND4 (N6016, N6011, N486, N848, N2100);
buf BUF1 (N6017, N6013);
nand NAND4 (N6018, N6016, N2587, N2110, N4558);
and AND3 (N6019, N6014, N2816, N540);
nor NOR4 (N6020, N5991, N5136, N3624, N4848);
or OR4 (N6021, N6018, N4163, N2361, N4014);
xor XOR2 (N6022, N6012, N3354);
xor XOR2 (N6023, N5998, N4919);
xor XOR2 (N6024, N6017, N3628);
buf BUF1 (N6025, N6006);
or OR3 (N6026, N6024, N1720, N3083);
or OR4 (N6027, N6020, N893, N4185, N3616);
and AND2 (N6028, N6008, N6005);
buf BUF1 (N6029, N5999);
and AND4 (N6030, N6019, N4244, N552, N2065);
nand NAND2 (N6031, N6029, N1692);
buf BUF1 (N6032, N6025);
or OR4 (N6033, N6032, N272, N5632, N5614);
and AND4 (N6034, N6033, N3214, N2809, N4513);
nand NAND4 (N6035, N6015, N114, N3980, N319);
buf BUF1 (N6036, N6022);
buf BUF1 (N6037, N6026);
buf BUF1 (N6038, N6035);
and AND4 (N6039, N6034, N3615, N1081, N5059);
not NOT1 (N6040, N6037);
nand NAND4 (N6041, N6030, N2823, N2185, N4844);
xor XOR2 (N6042, N6031, N2205);
nor NOR4 (N6043, N6039, N1446, N1913, N3411);
and AND3 (N6044, N6041, N4019, N1375);
not NOT1 (N6045, N6042);
xor XOR2 (N6046, N6023, N1093);
not NOT1 (N6047, N6043);
not NOT1 (N6048, N6044);
and AND3 (N6049, N6021, N3112, N2325);
nand NAND4 (N6050, N6049, N5247, N284, N5252);
and AND2 (N6051, N6046, N2166);
buf BUF1 (N6052, N6050);
buf BUF1 (N6053, N6040);
not NOT1 (N6054, N6028);
nand NAND2 (N6055, N6047, N4887);
nor NOR2 (N6056, N6051, N2560);
not NOT1 (N6057, N6053);
xor XOR2 (N6058, N6036, N1966);
or OR4 (N6059, N6058, N2104, N5935, N1804);
and AND2 (N6060, N6056, N4963);
nor NOR4 (N6061, N6060, N3294, N3729, N4466);
xor XOR2 (N6062, N6027, N179);
nand NAND4 (N6063, N6038, N2770, N1716, N4412);
xor XOR2 (N6064, N6057, N2485);
nand NAND4 (N6065, N6059, N397, N768, N3617);
nor NOR4 (N6066, N6061, N4934, N4626, N5970);
nor NOR2 (N6067, N6045, N5092);
buf BUF1 (N6068, N6063);
not NOT1 (N6069, N6066);
and AND4 (N6070, N6054, N728, N1549, N4162);
and AND4 (N6071, N6064, N2933, N4093, N393);
or OR2 (N6072, N6068, N3419);
buf BUF1 (N6073, N6070);
nand NAND3 (N6074, N6067, N3353, N4376);
nor NOR2 (N6075, N6069, N1464);
and AND3 (N6076, N6071, N2662, N4269);
buf BUF1 (N6077, N6073);
nor NOR2 (N6078, N6048, N253);
xor XOR2 (N6079, N6075, N1583);
buf BUF1 (N6080, N6055);
nand NAND3 (N6081, N6074, N4014, N3752);
nor NOR4 (N6082, N6079, N2072, N3813, N4011);
buf BUF1 (N6083, N6081);
nor NOR3 (N6084, N6062, N477, N3759);
nor NOR4 (N6085, N6076, N1239, N5223, N3274);
xor XOR2 (N6086, N6084, N4814);
nor NOR4 (N6087, N6082, N4518, N663, N4594);
or OR3 (N6088, N6085, N3160, N1526);
nand NAND2 (N6089, N6052, N3353);
nand NAND2 (N6090, N6088, N3709);
nand NAND4 (N6091, N6090, N4332, N1918, N2233);
or OR2 (N6092, N6077, N1412);
and AND3 (N6093, N6080, N2641, N3625);
xor XOR2 (N6094, N6078, N1087);
and AND3 (N6095, N6072, N391, N4750);
and AND2 (N6096, N6092, N4822);
or OR3 (N6097, N6089, N1495, N1077);
nand NAND3 (N6098, N6091, N5817, N461);
buf BUF1 (N6099, N6097);
not NOT1 (N6100, N6087);
or OR2 (N6101, N6086, N2526);
nand NAND2 (N6102, N6083, N2909);
nor NOR2 (N6103, N6093, N5089);
and AND4 (N6104, N6098, N4296, N4245, N2348);
not NOT1 (N6105, N6099);
not NOT1 (N6106, N6095);
nor NOR2 (N6107, N6100, N3732);
and AND4 (N6108, N6103, N2501, N893, N4660);
nor NOR4 (N6109, N6101, N2184, N412, N4391);
and AND3 (N6110, N6107, N5150, N2823);
nor NOR2 (N6111, N6104, N2534);
or OR4 (N6112, N6065, N5089, N5600, N63);
and AND2 (N6113, N6105, N2533);
not NOT1 (N6114, N6110);
not NOT1 (N6115, N6108);
and AND3 (N6116, N6115, N2401, N5916);
nor NOR3 (N6117, N6106, N1584, N560);
xor XOR2 (N6118, N6094, N2812);
xor XOR2 (N6119, N6109, N3057);
not NOT1 (N6120, N6117);
nand NAND4 (N6121, N6116, N770, N1340, N1686);
buf BUF1 (N6122, N6121);
xor XOR2 (N6123, N6112, N2990);
nor NOR2 (N6124, N6119, N5047);
xor XOR2 (N6125, N6124, N183);
nand NAND2 (N6126, N6123, N872);
nor NOR3 (N6127, N6125, N4841, N1376);
or OR3 (N6128, N6114, N1370, N1907);
nor NOR4 (N6129, N6128, N1839, N2956, N3304);
xor XOR2 (N6130, N6126, N293);
and AND4 (N6131, N6118, N584, N1802, N3992);
nor NOR3 (N6132, N6130, N4245, N4548);
xor XOR2 (N6133, N6102, N2388);
and AND4 (N6134, N6111, N4896, N5083, N1413);
or OR2 (N6135, N6131, N5899);
and AND3 (N6136, N6129, N6050, N2298);
not NOT1 (N6137, N6122);
xor XOR2 (N6138, N6096, N3283);
not NOT1 (N6139, N6132);
nand NAND4 (N6140, N6134, N4346, N2591, N5986);
not NOT1 (N6141, N6113);
buf BUF1 (N6142, N6140);
nand NAND4 (N6143, N6142, N1156, N2311, N4928);
not NOT1 (N6144, N6120);
nand NAND3 (N6145, N6138, N5815, N3414);
buf BUF1 (N6146, N6133);
buf BUF1 (N6147, N6145);
nor NOR4 (N6148, N6136, N1145, N563, N452);
not NOT1 (N6149, N6148);
nor NOR3 (N6150, N6127, N92, N4898);
and AND3 (N6151, N6135, N1222, N2830);
buf BUF1 (N6152, N6141);
not NOT1 (N6153, N6151);
nand NAND2 (N6154, N6146, N1066);
buf BUF1 (N6155, N6153);
and AND3 (N6156, N6139, N2130, N4608);
buf BUF1 (N6157, N6155);
xor XOR2 (N6158, N6157, N1724);
or OR2 (N6159, N6150, N3695);
xor XOR2 (N6160, N6147, N2285);
and AND4 (N6161, N6160, N3467, N1972, N5000);
xor XOR2 (N6162, N6158, N1303);
or OR2 (N6163, N6159, N2153);
not NOT1 (N6164, N6152);
xor XOR2 (N6165, N6143, N793);
and AND3 (N6166, N6154, N4957, N5454);
and AND3 (N6167, N6164, N5871, N2482);
nand NAND4 (N6168, N6137, N5285, N2797, N3899);
and AND2 (N6169, N6168, N2796);
xor XOR2 (N6170, N6144, N75);
nand NAND2 (N6171, N6170, N6039);
or OR3 (N6172, N6161, N5453, N4559);
nor NOR2 (N6173, N6167, N1513);
nand NAND4 (N6174, N6156, N4225, N3510, N2702);
xor XOR2 (N6175, N6165, N1366);
and AND4 (N6176, N6149, N1830, N5029, N2651);
and AND2 (N6177, N6173, N6099);
xor XOR2 (N6178, N6166, N3448);
not NOT1 (N6179, N6171);
xor XOR2 (N6180, N6177, N3890);
buf BUF1 (N6181, N6174);
buf BUF1 (N6182, N6181);
buf BUF1 (N6183, N6169);
nor NOR3 (N6184, N6180, N3780, N2785);
buf BUF1 (N6185, N6182);
nand NAND2 (N6186, N6185, N4505);
or OR2 (N6187, N6183, N2649);
nor NOR4 (N6188, N6178, N1629, N1030, N2918);
xor XOR2 (N6189, N6175, N6);
nor NOR3 (N6190, N6163, N5206, N2358);
nand NAND2 (N6191, N6172, N4766);
not NOT1 (N6192, N6191);
nor NOR3 (N6193, N6189, N383, N6065);
and AND3 (N6194, N6179, N36, N5349);
or OR4 (N6195, N6194, N5315, N3723, N4644);
and AND3 (N6196, N6192, N140, N4170);
nor NOR2 (N6197, N6195, N539);
or OR4 (N6198, N6162, N1357, N4071, N3627);
buf BUF1 (N6199, N6198);
nand NAND2 (N6200, N6176, N1048);
and AND3 (N6201, N6193, N2788, N5403);
buf BUF1 (N6202, N6186);
buf BUF1 (N6203, N6202);
and AND2 (N6204, N6188, N574);
nor NOR4 (N6205, N6203, N2538, N5636, N3278);
buf BUF1 (N6206, N6201);
buf BUF1 (N6207, N6184);
xor XOR2 (N6208, N6200, N3273);
xor XOR2 (N6209, N6199, N4840);
or OR4 (N6210, N6209, N1448, N2192, N6122);
and AND2 (N6211, N6206, N656);
xor XOR2 (N6212, N6210, N4943);
nor NOR4 (N6213, N6212, N5645, N6019, N1173);
or OR4 (N6214, N6211, N2496, N2255, N2465);
buf BUF1 (N6215, N6213);
nor NOR3 (N6216, N6204, N3170, N3994);
nand NAND2 (N6217, N6214, N5858);
xor XOR2 (N6218, N6190, N275);
nand NAND4 (N6219, N6216, N2952, N4673, N2326);
buf BUF1 (N6220, N6215);
and AND2 (N6221, N6207, N4929);
not NOT1 (N6222, N6208);
nor NOR3 (N6223, N6219, N4619, N5175);
buf BUF1 (N6224, N6223);
nand NAND3 (N6225, N6187, N101, N5200);
not NOT1 (N6226, N6197);
or OR2 (N6227, N6222, N4711);
nor NOR2 (N6228, N6196, N5497);
buf BUF1 (N6229, N6226);
nor NOR3 (N6230, N6225, N2060, N4753);
and AND3 (N6231, N6220, N5182, N3944);
nand NAND2 (N6232, N6230, N3082);
or OR2 (N6233, N6229, N4743);
xor XOR2 (N6234, N6232, N4338);
nand NAND3 (N6235, N6231, N2159, N3734);
not NOT1 (N6236, N6234);
not NOT1 (N6237, N6217);
nor NOR2 (N6238, N6218, N5091);
nand NAND4 (N6239, N6237, N2942, N272, N5528);
nor NOR3 (N6240, N6228, N4490, N5666);
or OR4 (N6241, N6221, N5850, N610, N5194);
not NOT1 (N6242, N6239);
xor XOR2 (N6243, N6224, N1608);
xor XOR2 (N6244, N6238, N812);
or OR4 (N6245, N6227, N5467, N4544, N2316);
nand NAND4 (N6246, N6245, N3753, N2782, N4686);
buf BUF1 (N6247, N6240);
buf BUF1 (N6248, N6242);
xor XOR2 (N6249, N6243, N3757);
nor NOR3 (N6250, N6247, N3755, N1597);
nor NOR4 (N6251, N6250, N2566, N1439, N345);
buf BUF1 (N6252, N6248);
and AND4 (N6253, N6249, N1451, N1131, N3025);
nor NOR2 (N6254, N6252, N1792);
and AND2 (N6255, N6251, N2610);
and AND4 (N6256, N6205, N3038, N4176, N2213);
nand NAND4 (N6257, N6253, N771, N3934, N2468);
nand NAND2 (N6258, N6244, N1848);
xor XOR2 (N6259, N6257, N2693);
nand NAND4 (N6260, N6246, N4378, N4989, N3132);
and AND4 (N6261, N6255, N5105, N1161, N4487);
or OR3 (N6262, N6260, N4963, N1361);
nand NAND4 (N6263, N6256, N4987, N4840, N736);
and AND2 (N6264, N6236, N4709);
nor NOR2 (N6265, N6264, N4551);
or OR4 (N6266, N6263, N1231, N476, N5046);
not NOT1 (N6267, N6254);
nor NOR2 (N6268, N6241, N2125);
or OR4 (N6269, N6235, N3527, N3083, N2623);
nand NAND2 (N6270, N6265, N1120);
nand NAND2 (N6271, N6269, N1209);
or OR2 (N6272, N6233, N4229);
not NOT1 (N6273, N6267);
or OR4 (N6274, N6261, N1895, N5313, N4377);
nand NAND4 (N6275, N6273, N4856, N4725, N2709);
buf BUF1 (N6276, N6268);
nor NOR3 (N6277, N6259, N3144, N1754);
xor XOR2 (N6278, N6266, N2895);
xor XOR2 (N6279, N6278, N4045);
xor XOR2 (N6280, N6277, N4443);
xor XOR2 (N6281, N6275, N3443);
or OR4 (N6282, N6274, N6260, N1005, N3163);
or OR4 (N6283, N6276, N4893, N351, N69);
nand NAND2 (N6284, N6283, N3077);
nand NAND4 (N6285, N6258, N543, N4327, N6155);
and AND4 (N6286, N6281, N5027, N2479, N3247);
not NOT1 (N6287, N6284);
and AND2 (N6288, N6270, N3229);
nor NOR4 (N6289, N6279, N1986, N312, N5137);
not NOT1 (N6290, N6282);
not NOT1 (N6291, N6272);
or OR2 (N6292, N6289, N1496);
and AND4 (N6293, N6292, N1757, N4403, N6167);
nand NAND4 (N6294, N6271, N2385, N2500, N3016);
xor XOR2 (N6295, N6293, N6033);
xor XOR2 (N6296, N6288, N5918);
and AND4 (N6297, N6295, N2514, N416, N5580);
buf BUF1 (N6298, N6297);
xor XOR2 (N6299, N6296, N4148);
xor XOR2 (N6300, N6262, N4173);
buf BUF1 (N6301, N6286);
and AND4 (N6302, N6298, N5262, N260, N2766);
not NOT1 (N6303, N6285);
not NOT1 (N6304, N6300);
or OR4 (N6305, N6291, N3949, N2194, N593);
nand NAND2 (N6306, N6301, N4007);
not NOT1 (N6307, N6299);
nand NAND3 (N6308, N6280, N6300, N1816);
nand NAND3 (N6309, N6304, N4190, N5493);
or OR3 (N6310, N6290, N795, N3424);
nand NAND4 (N6311, N6306, N2592, N1562, N1427);
xor XOR2 (N6312, N6287, N4876);
nand NAND2 (N6313, N6311, N1871);
or OR3 (N6314, N6307, N2513, N2895);
and AND3 (N6315, N6309, N2695, N5686);
not NOT1 (N6316, N6314);
buf BUF1 (N6317, N6313);
nand NAND4 (N6318, N6315, N805, N2835, N5973);
or OR2 (N6319, N6318, N50);
xor XOR2 (N6320, N6317, N4162);
xor XOR2 (N6321, N6302, N1364);
not NOT1 (N6322, N6312);
or OR4 (N6323, N6316, N1469, N1533, N5350);
xor XOR2 (N6324, N6320, N2877);
nor NOR3 (N6325, N6310, N3135, N3634);
nor NOR2 (N6326, N6303, N3590);
xor XOR2 (N6327, N6323, N39);
nand NAND3 (N6328, N6308, N5298, N4521);
nand NAND3 (N6329, N6325, N591, N1825);
or OR2 (N6330, N6326, N1104);
nand NAND4 (N6331, N6324, N5842, N252, N4410);
nor NOR2 (N6332, N6331, N6306);
nand NAND4 (N6333, N6332, N5223, N5361, N1873);
not NOT1 (N6334, N6333);
nor NOR4 (N6335, N6322, N5160, N3109, N5561);
buf BUF1 (N6336, N6294);
nor NOR2 (N6337, N6330, N872);
and AND4 (N6338, N6334, N185, N5904, N1288);
not NOT1 (N6339, N6335);
xor XOR2 (N6340, N6329, N1741);
nand NAND4 (N6341, N6328, N950, N1941, N3913);
buf BUF1 (N6342, N6319);
and AND2 (N6343, N6340, N815);
not NOT1 (N6344, N6342);
nand NAND2 (N6345, N6305, N5567);
not NOT1 (N6346, N6345);
nand NAND2 (N6347, N6321, N3316);
or OR2 (N6348, N6346, N732);
buf BUF1 (N6349, N6344);
nand NAND3 (N6350, N6327, N594, N86);
nor NOR3 (N6351, N6349, N5145, N2747);
nand NAND3 (N6352, N6336, N4211, N2551);
nand NAND4 (N6353, N6348, N73, N2777, N5713);
buf BUF1 (N6354, N6339);
buf BUF1 (N6355, N6338);
buf BUF1 (N6356, N6341);
or OR3 (N6357, N6337, N5715, N1098);
not NOT1 (N6358, N6350);
xor XOR2 (N6359, N6353, N1907);
not NOT1 (N6360, N6343);
or OR4 (N6361, N6352, N3576, N5335, N2075);
not NOT1 (N6362, N6354);
not NOT1 (N6363, N6347);
nand NAND2 (N6364, N6360, N2401);
nand NAND4 (N6365, N6364, N3625, N4451, N3121);
not NOT1 (N6366, N6365);
not NOT1 (N6367, N6356);
nand NAND4 (N6368, N6366, N3910, N1696, N4721);
and AND4 (N6369, N6359, N6332, N5141, N4060);
or OR2 (N6370, N6351, N5046);
nor NOR2 (N6371, N6362, N177);
nand NAND3 (N6372, N6370, N4097, N6349);
or OR4 (N6373, N6369, N1643, N1731, N166);
nor NOR4 (N6374, N6373, N2063, N430, N4899);
nand NAND2 (N6375, N6357, N2502);
or OR3 (N6376, N6374, N599, N2819);
nor NOR2 (N6377, N6355, N846);
xor XOR2 (N6378, N6372, N2793);
nor NOR2 (N6379, N6376, N5008);
xor XOR2 (N6380, N6363, N3483);
not NOT1 (N6381, N6367);
and AND4 (N6382, N6375, N1411, N448, N850);
nor NOR2 (N6383, N6382, N5135);
not NOT1 (N6384, N6383);
xor XOR2 (N6385, N6358, N2523);
not NOT1 (N6386, N6384);
nor NOR4 (N6387, N6380, N3223, N3938, N5189);
or OR4 (N6388, N6361, N6332, N2581, N5158);
not NOT1 (N6389, N6381);
xor XOR2 (N6390, N6389, N2897);
not NOT1 (N6391, N6385);
buf BUF1 (N6392, N6368);
nand NAND2 (N6393, N6379, N5637);
buf BUF1 (N6394, N6393);
not NOT1 (N6395, N6377);
buf BUF1 (N6396, N6386);
or OR4 (N6397, N6395, N3833, N3298, N3883);
not NOT1 (N6398, N6371);
buf BUF1 (N6399, N6391);
or OR2 (N6400, N6398, N5154);
nand NAND2 (N6401, N6390, N4949);
xor XOR2 (N6402, N6399, N4174);
not NOT1 (N6403, N6394);
nor NOR2 (N6404, N6403, N628);
nor NOR3 (N6405, N6378, N3514, N3511);
and AND4 (N6406, N6402, N1863, N4950, N2995);
buf BUF1 (N6407, N6397);
and AND4 (N6408, N6392, N807, N5125, N2868);
or OR4 (N6409, N6396, N3680, N3211, N5335);
or OR4 (N6410, N6405, N5317, N986, N4763);
or OR2 (N6411, N6404, N420);
nor NOR3 (N6412, N6407, N3609, N2358);
or OR2 (N6413, N6412, N4669);
not NOT1 (N6414, N6387);
xor XOR2 (N6415, N6408, N1993);
buf BUF1 (N6416, N6400);
xor XOR2 (N6417, N6388, N3036);
buf BUF1 (N6418, N6411);
nor NOR3 (N6419, N6406, N4758, N5133);
xor XOR2 (N6420, N6416, N5418);
xor XOR2 (N6421, N6401, N6237);
or OR4 (N6422, N6420, N4696, N426, N5709);
nand NAND3 (N6423, N6418, N1569, N3437);
not NOT1 (N6424, N6417);
nand NAND4 (N6425, N6424, N4272, N3231, N2150);
xor XOR2 (N6426, N6413, N2681);
nand NAND2 (N6427, N6409, N45);
nand NAND4 (N6428, N6415, N3218, N4704, N6258);
buf BUF1 (N6429, N6428);
buf BUF1 (N6430, N6419);
nand NAND3 (N6431, N6429, N3221, N810);
xor XOR2 (N6432, N6421, N2235);
nor NOR3 (N6433, N6425, N1224, N3837);
not NOT1 (N6434, N6432);
xor XOR2 (N6435, N6426, N1751);
and AND2 (N6436, N6431, N335);
or OR2 (N6437, N6436, N2792);
buf BUF1 (N6438, N6414);
buf BUF1 (N6439, N6423);
xor XOR2 (N6440, N6434, N3540);
buf BUF1 (N6441, N6439);
or OR3 (N6442, N6410, N2911, N2015);
nand NAND4 (N6443, N6438, N6276, N2757, N5);
and AND4 (N6444, N6430, N5169, N3099, N393);
or OR3 (N6445, N6437, N1131, N5232);
not NOT1 (N6446, N6444);
nor NOR4 (N6447, N6440, N2377, N5706, N5529);
nand NAND2 (N6448, N6435, N2531);
xor XOR2 (N6449, N6446, N1984);
or OR2 (N6450, N6441, N4606);
and AND4 (N6451, N6433, N959, N2462, N4640);
nand NAND3 (N6452, N6445, N3791, N6212);
or OR3 (N6453, N6451, N4697, N1326);
or OR2 (N6454, N6449, N3927);
not NOT1 (N6455, N6453);
xor XOR2 (N6456, N6450, N6333);
nand NAND2 (N6457, N6427, N4380);
or OR2 (N6458, N6448, N2167);
not NOT1 (N6459, N6442);
nor NOR3 (N6460, N6458, N1608, N2455);
buf BUF1 (N6461, N6454);
xor XOR2 (N6462, N6461, N6363);
and AND3 (N6463, N6447, N2639, N6345);
nor NOR4 (N6464, N6455, N1468, N1624, N1977);
and AND3 (N6465, N6457, N6371, N3451);
buf BUF1 (N6466, N6443);
nand NAND2 (N6467, N6463, N714);
nand NAND2 (N6468, N6452, N4241);
nand NAND4 (N6469, N6459, N971, N4809, N494);
xor XOR2 (N6470, N6468, N5957);
not NOT1 (N6471, N6465);
and AND4 (N6472, N6464, N960, N2043, N390);
buf BUF1 (N6473, N6462);
nand NAND2 (N6474, N6472, N71);
nand NAND3 (N6475, N6467, N2664, N2824);
nor NOR3 (N6476, N6469, N3857, N3367);
nand NAND2 (N6477, N6422, N4731);
nand NAND4 (N6478, N6460, N2116, N933, N808);
and AND4 (N6479, N6475, N4070, N5433, N3890);
not NOT1 (N6480, N6471);
not NOT1 (N6481, N6479);
buf BUF1 (N6482, N6478);
not NOT1 (N6483, N6466);
or OR4 (N6484, N6477, N4096, N4627, N346);
nand NAND3 (N6485, N6470, N1477, N4163);
nor NOR3 (N6486, N6456, N4499, N5480);
nand NAND4 (N6487, N6486, N2003, N937, N2047);
nand NAND3 (N6488, N6484, N1685, N2914);
not NOT1 (N6489, N6480);
not NOT1 (N6490, N6487);
buf BUF1 (N6491, N6482);
buf BUF1 (N6492, N6490);
buf BUF1 (N6493, N6481);
buf BUF1 (N6494, N6485);
or OR3 (N6495, N6489, N4151, N410);
and AND4 (N6496, N6494, N5327, N2145, N1139);
nor NOR3 (N6497, N6488, N749, N983);
buf BUF1 (N6498, N6497);
not NOT1 (N6499, N6473);
or OR2 (N6500, N6483, N6120);
not NOT1 (N6501, N6495);
and AND3 (N6502, N6492, N5579, N2469);
or OR2 (N6503, N6476, N3261);
buf BUF1 (N6504, N6499);
nand NAND3 (N6505, N6502, N1587, N6197);
xor XOR2 (N6506, N6493, N369);
nor NOR3 (N6507, N6500, N6493, N5237);
nor NOR3 (N6508, N6506, N5349, N4359);
buf BUF1 (N6509, N6496);
not NOT1 (N6510, N6491);
not NOT1 (N6511, N6507);
nand NAND2 (N6512, N6508, N4677);
or OR4 (N6513, N6474, N3875, N166, N3766);
xor XOR2 (N6514, N6510, N450);
nor NOR3 (N6515, N6505, N5330, N3997);
buf BUF1 (N6516, N6501);
buf BUF1 (N6517, N6509);
and AND3 (N6518, N6498, N3202, N1914);
xor XOR2 (N6519, N6504, N2353);
xor XOR2 (N6520, N6513, N1449);
xor XOR2 (N6521, N6520, N2773);
buf BUF1 (N6522, N6514);
nor NOR4 (N6523, N6516, N6338, N5350, N5335);
not NOT1 (N6524, N6522);
not NOT1 (N6525, N6518);
buf BUF1 (N6526, N6503);
buf BUF1 (N6527, N6525);
nand NAND3 (N6528, N6515, N315, N3977);
and AND3 (N6529, N6511, N3817, N4690);
and AND3 (N6530, N6526, N912, N2199);
nor NOR3 (N6531, N6530, N2838, N6126);
not NOT1 (N6532, N6523);
and AND3 (N6533, N6519, N3808, N1143);
nand NAND2 (N6534, N6528, N3342);
or OR4 (N6535, N6521, N5479, N5651, N332);
buf BUF1 (N6536, N6532);
not NOT1 (N6537, N6529);
and AND3 (N6538, N6534, N5616, N155);
not NOT1 (N6539, N6531);
nand NAND4 (N6540, N6527, N2837, N6510, N4902);
buf BUF1 (N6541, N6538);
nor NOR2 (N6542, N6536, N6044);
buf BUF1 (N6543, N6541);
not NOT1 (N6544, N6535);
xor XOR2 (N6545, N6544, N5042);
nor NOR4 (N6546, N6512, N2264, N571, N5360);
nor NOR4 (N6547, N6543, N3419, N5614, N5060);
nor NOR4 (N6548, N6540, N6249, N6327, N4267);
and AND2 (N6549, N6546, N6375);
nand NAND4 (N6550, N6542, N637, N3904, N4378);
nor NOR2 (N6551, N6547, N3769);
nor NOR4 (N6552, N6545, N4749, N1181, N6184);
nand NAND2 (N6553, N6549, N763);
buf BUF1 (N6554, N6524);
or OR3 (N6555, N6553, N5966, N4306);
xor XOR2 (N6556, N6539, N4231);
nand NAND2 (N6557, N6537, N384);
buf BUF1 (N6558, N6517);
nand NAND3 (N6559, N6555, N3804, N3830);
buf BUF1 (N6560, N6556);
nand NAND3 (N6561, N6552, N6461, N1174);
nand NAND3 (N6562, N6554, N97, N5788);
and AND4 (N6563, N6562, N3332, N4514, N3153);
or OR2 (N6564, N6559, N6170);
not NOT1 (N6565, N6560);
or OR3 (N6566, N6550, N4001, N1058);
nand NAND2 (N6567, N6565, N3343);
xor XOR2 (N6568, N6561, N2856);
buf BUF1 (N6569, N6548);
buf BUF1 (N6570, N6568);
not NOT1 (N6571, N6569);
not NOT1 (N6572, N6570);
xor XOR2 (N6573, N6551, N3138);
and AND2 (N6574, N6564, N1093);
not NOT1 (N6575, N6566);
nand NAND2 (N6576, N6574, N1397);
not NOT1 (N6577, N6576);
xor XOR2 (N6578, N6575, N428);
buf BUF1 (N6579, N6558);
nor NOR2 (N6580, N6567, N1367);
or OR4 (N6581, N6533, N1723, N2077, N6188);
and AND3 (N6582, N6580, N4408, N1140);
and AND4 (N6583, N6578, N606, N2921, N6017);
xor XOR2 (N6584, N6582, N3229);
nand NAND2 (N6585, N6584, N1577);
xor XOR2 (N6586, N6579, N559);
not NOT1 (N6587, N6563);
and AND3 (N6588, N6577, N2866, N564);
xor XOR2 (N6589, N6572, N4116);
xor XOR2 (N6590, N6588, N4689);
not NOT1 (N6591, N6585);
nand NAND3 (N6592, N6573, N3219, N673);
not NOT1 (N6593, N6586);
nand NAND4 (N6594, N6592, N2045, N2439, N3985);
xor XOR2 (N6595, N6587, N2467);
nand NAND2 (N6596, N6589, N790);
and AND3 (N6597, N6595, N4914, N2262);
xor XOR2 (N6598, N6594, N2515);
buf BUF1 (N6599, N6593);
buf BUF1 (N6600, N6581);
xor XOR2 (N6601, N6591, N3295);
buf BUF1 (N6602, N6597);
nand NAND2 (N6603, N6590, N2545);
nor NOR4 (N6604, N6598, N4729, N880, N3589);
or OR3 (N6605, N6600, N1687, N3655);
buf BUF1 (N6606, N6601);
nand NAND4 (N6607, N6599, N414, N1435, N448);
nor NOR3 (N6608, N6596, N3994, N5243);
or OR3 (N6609, N6604, N3400, N493);
nor NOR3 (N6610, N6571, N253, N4388);
nand NAND2 (N6611, N6557, N245);
and AND3 (N6612, N6607, N7, N1465);
buf BUF1 (N6613, N6603);
or OR2 (N6614, N6608, N4093);
nand NAND4 (N6615, N6583, N2815, N4066, N6512);
not NOT1 (N6616, N6606);
and AND2 (N6617, N6610, N2289);
xor XOR2 (N6618, N6613, N6265);
and AND3 (N6619, N6609, N167, N4814);
xor XOR2 (N6620, N6615, N5776);
nor NOR3 (N6621, N6618, N2621, N5872);
and AND3 (N6622, N6619, N1628, N6424);
or OR3 (N6623, N6620, N6172, N965);
and AND3 (N6624, N6621, N1714, N3346);
nor NOR3 (N6625, N6617, N4122, N5007);
not NOT1 (N6626, N6623);
or OR2 (N6627, N6612, N2557);
not NOT1 (N6628, N6616);
buf BUF1 (N6629, N6605);
buf BUF1 (N6630, N6611);
nand NAND3 (N6631, N6626, N5773, N1165);
or OR4 (N6632, N6627, N1839, N4832, N406);
or OR2 (N6633, N6629, N4727);
not NOT1 (N6634, N6631);
buf BUF1 (N6635, N6602);
not NOT1 (N6636, N6622);
nand NAND4 (N6637, N6624, N4364, N2529, N3685);
nand NAND3 (N6638, N6633, N2675, N4062);
nand NAND3 (N6639, N6638, N4654, N5623);
not NOT1 (N6640, N6636);
nor NOR3 (N6641, N6632, N181, N4678);
nand NAND4 (N6642, N6639, N1552, N3196, N3148);
nand NAND4 (N6643, N6635, N4194, N3320, N1396);
nor NOR4 (N6644, N6642, N5632, N1804, N2311);
not NOT1 (N6645, N6641);
nor NOR2 (N6646, N6643, N1243);
nand NAND4 (N6647, N6628, N5527, N3226, N702);
nor NOR4 (N6648, N6614, N998, N6153, N2655);
and AND2 (N6649, N6645, N3260);
nor NOR2 (N6650, N6647, N169);
nand NAND2 (N6651, N6640, N376);
buf BUF1 (N6652, N6637);
nor NOR2 (N6653, N6630, N1672);
not NOT1 (N6654, N6649);
buf BUF1 (N6655, N6650);
nor NOR4 (N6656, N6648, N2496, N760, N1448);
nor NOR4 (N6657, N6652, N1152, N5575, N4923);
not NOT1 (N6658, N6625);
xor XOR2 (N6659, N6646, N6074);
or OR3 (N6660, N6657, N2038, N5015);
xor XOR2 (N6661, N6655, N4789);
not NOT1 (N6662, N6654);
and AND4 (N6663, N6644, N3207, N5161, N2376);
and AND3 (N6664, N6660, N2799, N2039);
or OR4 (N6665, N6656, N2528, N5925, N1620);
buf BUF1 (N6666, N6659);
buf BUF1 (N6667, N6653);
xor XOR2 (N6668, N6661, N3575);
nor NOR3 (N6669, N6651, N5336, N1869);
nor NOR2 (N6670, N6666, N884);
nor NOR3 (N6671, N6663, N5102, N481);
nor NOR3 (N6672, N6667, N238, N965);
nand NAND2 (N6673, N6658, N3842);
not NOT1 (N6674, N6668);
nand NAND4 (N6675, N6665, N5260, N3836, N6512);
nor NOR2 (N6676, N6675, N1435);
not NOT1 (N6677, N6634);
buf BUF1 (N6678, N6662);
nor NOR3 (N6679, N6669, N6365, N2298);
or OR2 (N6680, N6679, N5440);
and AND3 (N6681, N6677, N6046, N5455);
and AND2 (N6682, N6676, N4673);
nand NAND4 (N6683, N6670, N4368, N4091, N3382);
buf BUF1 (N6684, N6664);
or OR3 (N6685, N6671, N3860, N262);
nor NOR2 (N6686, N6674, N591);
nor NOR2 (N6687, N6683, N52);
or OR4 (N6688, N6672, N4169, N5968, N534);
buf BUF1 (N6689, N6682);
buf BUF1 (N6690, N6680);
nor NOR4 (N6691, N6686, N1044, N930, N1449);
nand NAND3 (N6692, N6684, N5030, N4529);
buf BUF1 (N6693, N6691);
nor NOR2 (N6694, N6681, N1501);
not NOT1 (N6695, N6689);
xor XOR2 (N6696, N6678, N5172);
nor NOR2 (N6697, N6687, N2537);
and AND4 (N6698, N6695, N2240, N802, N40);
not NOT1 (N6699, N6693);
nor NOR4 (N6700, N6698, N28, N5388, N4423);
xor XOR2 (N6701, N6692, N2827);
nand NAND2 (N6702, N6697, N3244);
xor XOR2 (N6703, N6700, N1824);
or OR3 (N6704, N6702, N1221, N6479);
buf BUF1 (N6705, N6694);
buf BUF1 (N6706, N6696);
and AND3 (N6707, N6706, N4325, N796);
not NOT1 (N6708, N6699);
nor NOR3 (N6709, N6705, N6426, N370);
nor NOR3 (N6710, N6690, N26, N5881);
nor NOR2 (N6711, N6704, N77);
and AND4 (N6712, N6685, N648, N1839, N310);
nor NOR4 (N6713, N6711, N6178, N2796, N2791);
xor XOR2 (N6714, N6688, N3798);
xor XOR2 (N6715, N6712, N2788);
buf BUF1 (N6716, N6703);
and AND3 (N6717, N6709, N4310, N3724);
buf BUF1 (N6718, N6708);
nor NOR4 (N6719, N6715, N3036, N6110, N188);
nor NOR2 (N6720, N6710, N3405);
and AND2 (N6721, N6717, N2164);
xor XOR2 (N6722, N6714, N1763);
and AND4 (N6723, N6722, N2045, N2459, N1607);
nand NAND2 (N6724, N6701, N4517);
buf BUF1 (N6725, N6713);
or OR2 (N6726, N6718, N4393);
and AND2 (N6727, N6726, N4758);
nor NOR4 (N6728, N6719, N4035, N5816, N1467);
and AND2 (N6729, N6721, N5632);
buf BUF1 (N6730, N6673);
or OR4 (N6731, N6716, N4855, N391, N3072);
buf BUF1 (N6732, N6707);
nand NAND3 (N6733, N6724, N2019, N3942);
xor XOR2 (N6734, N6728, N5872);
or OR4 (N6735, N6725, N1704, N1479, N5903);
and AND4 (N6736, N6732, N5787, N6232, N4412);
buf BUF1 (N6737, N6723);
or OR3 (N6738, N6735, N1951, N374);
nand NAND2 (N6739, N6733, N2179);
nor NOR4 (N6740, N6731, N2498, N4556, N1629);
and AND4 (N6741, N6730, N5932, N5195, N1094);
nand NAND2 (N6742, N6727, N6181);
not NOT1 (N6743, N6738);
xor XOR2 (N6744, N6720, N3605);
and AND3 (N6745, N6742, N4547, N4167);
or OR4 (N6746, N6745, N4400, N5847, N5494);
not NOT1 (N6747, N6744);
and AND4 (N6748, N6746, N1953, N4325, N5939);
and AND3 (N6749, N6729, N5205, N5818);
and AND3 (N6750, N6739, N4968, N3478);
buf BUF1 (N6751, N6749);
or OR2 (N6752, N6736, N5226);
or OR3 (N6753, N6752, N3881, N958);
not NOT1 (N6754, N6741);
xor XOR2 (N6755, N6753, N183);
and AND4 (N6756, N6754, N3864, N1578, N3920);
not NOT1 (N6757, N6751);
xor XOR2 (N6758, N6740, N5849);
nor NOR3 (N6759, N6756, N2193, N2002);
xor XOR2 (N6760, N6750, N969);
not NOT1 (N6761, N6734);
or OR2 (N6762, N6761, N888);
or OR3 (N6763, N6758, N3959, N3963);
and AND4 (N6764, N6737, N828, N9, N369);
not NOT1 (N6765, N6755);
not NOT1 (N6766, N6759);
not NOT1 (N6767, N6766);
nor NOR4 (N6768, N6747, N71, N3536, N2245);
nor NOR2 (N6769, N6743, N2569);
and AND3 (N6770, N6748, N3708, N3953);
and AND2 (N6771, N6769, N1234);
nor NOR4 (N6772, N6770, N4381, N4706, N3457);
nand NAND2 (N6773, N6767, N1956);
not NOT1 (N6774, N6760);
not NOT1 (N6775, N6768);
and AND4 (N6776, N6765, N415, N2421, N391);
or OR3 (N6777, N6757, N3423, N3942);
or OR3 (N6778, N6763, N3679, N6094);
xor XOR2 (N6779, N6776, N1857);
nand NAND3 (N6780, N6773, N3016, N6486);
nand NAND4 (N6781, N6762, N1901, N3384, N3969);
or OR4 (N6782, N6771, N2959, N6438, N3135);
not NOT1 (N6783, N6780);
and AND4 (N6784, N6772, N6198, N4918, N5592);
nor NOR3 (N6785, N6764, N3653, N1010);
buf BUF1 (N6786, N6781);
or OR4 (N6787, N6782, N659, N6531, N3628);
not NOT1 (N6788, N6786);
not NOT1 (N6789, N6778);
buf BUF1 (N6790, N6779);
buf BUF1 (N6791, N6788);
not NOT1 (N6792, N6789);
xor XOR2 (N6793, N6784, N5429);
nand NAND3 (N6794, N6785, N5450, N3049);
not NOT1 (N6795, N6777);
and AND4 (N6796, N6793, N279, N3196, N1472);
not NOT1 (N6797, N6774);
buf BUF1 (N6798, N6794);
buf BUF1 (N6799, N6783);
buf BUF1 (N6800, N6796);
xor XOR2 (N6801, N6798, N5964);
xor XOR2 (N6802, N6792, N5951);
buf BUF1 (N6803, N6795);
buf BUF1 (N6804, N6803);
not NOT1 (N6805, N6791);
not NOT1 (N6806, N6790);
nor NOR4 (N6807, N6806, N6508, N4395, N1805);
or OR2 (N6808, N6807, N1109);
or OR2 (N6809, N6775, N3737);
buf BUF1 (N6810, N6801);
nor NOR4 (N6811, N6809, N2561, N35, N5366);
nor NOR2 (N6812, N6800, N4227);
or OR3 (N6813, N6804, N1720, N347);
xor XOR2 (N6814, N6811, N4971);
buf BUF1 (N6815, N6808);
not NOT1 (N6816, N6805);
xor XOR2 (N6817, N6815, N6601);
xor XOR2 (N6818, N6817, N6340);
xor XOR2 (N6819, N6816, N3928);
and AND4 (N6820, N6787, N1534, N6192, N506);
nor NOR3 (N6821, N6797, N1681, N6501);
or OR2 (N6822, N6819, N1935);
buf BUF1 (N6823, N6822);
xor XOR2 (N6824, N6814, N2372);
or OR4 (N6825, N6820, N1485, N1750, N2651);
not NOT1 (N6826, N6818);
xor XOR2 (N6827, N6802, N1396);
xor XOR2 (N6828, N6827, N467);
or OR2 (N6829, N6821, N2779);
nand NAND4 (N6830, N6826, N2437, N5986, N3913);
and AND3 (N6831, N6823, N1519, N4429);
xor XOR2 (N6832, N6830, N257);
nor NOR4 (N6833, N6825, N4681, N4205, N236);
or OR2 (N6834, N6833, N2058);
and AND2 (N6835, N6799, N5552);
nor NOR3 (N6836, N6832, N6416, N4592);
and AND4 (N6837, N6831, N1270, N3505, N3428);
or OR3 (N6838, N6828, N161, N78);
nor NOR2 (N6839, N6837, N1294);
buf BUF1 (N6840, N6824);
nand NAND2 (N6841, N6839, N2880);
nor NOR3 (N6842, N6812, N5547, N856);
and AND3 (N6843, N6810, N2650, N6401);
or OR3 (N6844, N6840, N1909, N3435);
or OR4 (N6845, N6841, N5014, N671, N980);
or OR3 (N6846, N6842, N1144, N4861);
nand NAND3 (N6847, N6844, N3857, N1027);
xor XOR2 (N6848, N6813, N1439);
not NOT1 (N6849, N6829);
or OR4 (N6850, N6849, N1253, N5215, N4828);
or OR4 (N6851, N6845, N4419, N5389, N5286);
buf BUF1 (N6852, N6835);
nand NAND3 (N6853, N6838, N6680, N1446);
nor NOR3 (N6854, N6843, N5322, N748);
nand NAND2 (N6855, N6836, N3815);
nor NOR4 (N6856, N6851, N4644, N2076, N4826);
xor XOR2 (N6857, N6855, N1552);
not NOT1 (N6858, N6850);
nor NOR2 (N6859, N6852, N1855);
buf BUF1 (N6860, N6853);
nor NOR3 (N6861, N6859, N2366, N822);
not NOT1 (N6862, N6860);
xor XOR2 (N6863, N6857, N671);
or OR4 (N6864, N6847, N3915, N3158, N3956);
nor NOR3 (N6865, N6856, N4438, N4527);
nand NAND2 (N6866, N6834, N6694);
buf BUF1 (N6867, N6848);
not NOT1 (N6868, N6866);
nor NOR4 (N6869, N6867, N5265, N3776, N5808);
xor XOR2 (N6870, N6854, N2839);
not NOT1 (N6871, N6865);
not NOT1 (N6872, N6870);
or OR4 (N6873, N6846, N1746, N4643, N4179);
buf BUF1 (N6874, N6873);
not NOT1 (N6875, N6869);
buf BUF1 (N6876, N6863);
buf BUF1 (N6877, N6874);
buf BUF1 (N6878, N6875);
or OR3 (N6879, N6861, N3826, N266);
nand NAND4 (N6880, N6876, N3328, N1526, N2742);
buf BUF1 (N6881, N6862);
xor XOR2 (N6882, N6879, N3850);
xor XOR2 (N6883, N6868, N3436);
xor XOR2 (N6884, N6883, N1839);
not NOT1 (N6885, N6884);
nor NOR4 (N6886, N6881, N2968, N442, N5074);
or OR4 (N6887, N6882, N3521, N2406, N5312);
or OR3 (N6888, N6877, N6098, N3982);
not NOT1 (N6889, N6887);
nor NOR3 (N6890, N6864, N5739, N6124);
not NOT1 (N6891, N6885);
buf BUF1 (N6892, N6889);
buf BUF1 (N6893, N6880);
or OR3 (N6894, N6890, N1827, N2592);
xor XOR2 (N6895, N6878, N5145);
and AND2 (N6896, N6891, N5846);
nor NOR2 (N6897, N6892, N263);
and AND4 (N6898, N6872, N3528, N5540, N3519);
or OR4 (N6899, N6895, N4415, N5811, N5292);
xor XOR2 (N6900, N6898, N5517);
nor NOR3 (N6901, N6871, N1819, N1572);
xor XOR2 (N6902, N6886, N3827);
or OR2 (N6903, N6901, N5862);
nor NOR4 (N6904, N6900, N4791, N3322, N4602);
buf BUF1 (N6905, N6897);
and AND2 (N6906, N6894, N3444);
nand NAND2 (N6907, N6893, N866);
nor NOR4 (N6908, N6896, N1465, N3614, N5488);
not NOT1 (N6909, N6908);
and AND4 (N6910, N6903, N5026, N5341, N2109);
or OR3 (N6911, N6899, N5381, N390);
nor NOR2 (N6912, N6909, N6270);
xor XOR2 (N6913, N6904, N3169);
not NOT1 (N6914, N6907);
nor NOR2 (N6915, N6906, N5318);
nor NOR3 (N6916, N6910, N1290, N5473);
nand NAND3 (N6917, N6888, N6195, N5254);
or OR2 (N6918, N6915, N5170);
xor XOR2 (N6919, N6911, N3425);
buf BUF1 (N6920, N6905);
nor NOR4 (N6921, N6918, N2038, N5677, N2719);
nand NAND3 (N6922, N6919, N214, N4934);
nand NAND4 (N6923, N6921, N4519, N5426, N3928);
buf BUF1 (N6924, N6916);
and AND2 (N6925, N6917, N3410);
nand NAND2 (N6926, N6924, N5902);
nor NOR4 (N6927, N6922, N826, N4236, N6631);
or OR2 (N6928, N6925, N6899);
xor XOR2 (N6929, N6912, N3172);
nand NAND2 (N6930, N6920, N1221);
xor XOR2 (N6931, N6923, N5658);
nand NAND4 (N6932, N6926, N1033, N6540, N871);
not NOT1 (N6933, N6902);
xor XOR2 (N6934, N6931, N5762);
nor NOR4 (N6935, N6914, N1942, N4260, N5335);
buf BUF1 (N6936, N6927);
or OR3 (N6937, N6858, N1862, N5608);
not NOT1 (N6938, N6934);
nand NAND4 (N6939, N6937, N1741, N4151, N5709);
xor XOR2 (N6940, N6935, N4314);
xor XOR2 (N6941, N6940, N3965);
and AND4 (N6942, N6938, N2835, N6103, N5324);
nor NOR4 (N6943, N6928, N5779, N1154, N115);
buf BUF1 (N6944, N6939);
xor XOR2 (N6945, N6929, N6004);
xor XOR2 (N6946, N6936, N3702);
nand NAND2 (N6947, N6945, N2007);
nand NAND2 (N6948, N6943, N2488);
buf BUF1 (N6949, N6946);
buf BUF1 (N6950, N6913);
xor XOR2 (N6951, N6933, N1368);
and AND4 (N6952, N6930, N3385, N6007, N3850);
xor XOR2 (N6953, N6949, N5169);
not NOT1 (N6954, N6950);
xor XOR2 (N6955, N6942, N4747);
nor NOR3 (N6956, N6952, N1535, N4235);
nand NAND3 (N6957, N6955, N1640, N4441);
xor XOR2 (N6958, N6954, N4500);
xor XOR2 (N6959, N6948, N2073);
xor XOR2 (N6960, N6951, N865);
not NOT1 (N6961, N6953);
not NOT1 (N6962, N6959);
buf BUF1 (N6963, N6956);
nand NAND2 (N6964, N6932, N5501);
and AND2 (N6965, N6964, N2904);
nand NAND4 (N6966, N6963, N3871, N4562, N1697);
nand NAND4 (N6967, N6966, N2279, N1481, N4541);
not NOT1 (N6968, N6944);
nand NAND2 (N6969, N6941, N4400);
not NOT1 (N6970, N6958);
buf BUF1 (N6971, N6962);
buf BUF1 (N6972, N6965);
buf BUF1 (N6973, N6970);
xor XOR2 (N6974, N6969, N2409);
not NOT1 (N6975, N6971);
nor NOR3 (N6976, N6975, N6533, N2879);
or OR4 (N6977, N6972, N3940, N4214, N1284);
nor NOR4 (N6978, N6968, N6685, N2683, N6363);
not NOT1 (N6979, N6960);
xor XOR2 (N6980, N6978, N1053);
nor NOR4 (N6981, N6967, N103, N4876, N4210);
nand NAND2 (N6982, N6981, N6409);
buf BUF1 (N6983, N6982);
or OR3 (N6984, N6961, N5510, N1423);
xor XOR2 (N6985, N6983, N1651);
nor NOR4 (N6986, N6979, N6580, N4058, N4107);
not NOT1 (N6987, N6974);
and AND4 (N6988, N6973, N3347, N3863, N5271);
nor NOR3 (N6989, N6947, N477, N1927);
nor NOR3 (N6990, N6988, N3358, N2286);
xor XOR2 (N6991, N6990, N374);
nor NOR4 (N6992, N6976, N14, N4761, N4213);
or OR2 (N6993, N6986, N5447);
or OR4 (N6994, N6992, N5591, N3788, N2622);
nand NAND4 (N6995, N6994, N5952, N1554, N3827);
buf BUF1 (N6996, N6977);
buf BUF1 (N6997, N6995);
buf BUF1 (N6998, N6989);
xor XOR2 (N6999, N6997, N2283);
buf BUF1 (N7000, N6987);
nand NAND4 (N7001, N6996, N2159, N2457, N4168);
xor XOR2 (N7002, N6998, N583);
not NOT1 (N7003, N6980);
nor NOR2 (N7004, N6991, N787);
not NOT1 (N7005, N6993);
not NOT1 (N7006, N7001);
nand NAND2 (N7007, N7003, N5963);
nand NAND3 (N7008, N7000, N4040, N1127);
nand NAND3 (N7009, N7008, N1082, N3892);
nand NAND2 (N7010, N7005, N3606);
or OR3 (N7011, N6985, N2237, N4049);
nor NOR2 (N7012, N7007, N5121);
nand NAND4 (N7013, N6999, N4308, N6140, N3568);
nor NOR4 (N7014, N6957, N5281, N3196, N4862);
or OR3 (N7015, N7009, N3443, N4156);
and AND3 (N7016, N7010, N5352, N5404);
buf BUF1 (N7017, N6984);
and AND4 (N7018, N7013, N2635, N4436, N1856);
and AND4 (N7019, N7012, N290, N1640, N3644);
or OR3 (N7020, N7017, N4438, N1520);
and AND2 (N7021, N7019, N6219);
nand NAND4 (N7022, N7021, N1220, N2620, N1555);
and AND3 (N7023, N7002, N771, N4968);
or OR4 (N7024, N7018, N4096, N713, N1059);
xor XOR2 (N7025, N7024, N1854);
buf BUF1 (N7026, N7025);
or OR2 (N7027, N7020, N3448);
xor XOR2 (N7028, N7015, N740);
not NOT1 (N7029, N7016);
nor NOR4 (N7030, N7027, N6065, N5553, N1689);
not NOT1 (N7031, N7006);
or OR2 (N7032, N7022, N6055);
buf BUF1 (N7033, N7011);
nand NAND3 (N7034, N7014, N890, N1648);
nor NOR3 (N7035, N7033, N6410, N3377);
and AND3 (N7036, N7029, N2341, N4454);
xor XOR2 (N7037, N7035, N648);
buf BUF1 (N7038, N7030);
not NOT1 (N7039, N7028);
nor NOR4 (N7040, N7004, N882, N6087, N6491);
buf BUF1 (N7041, N7026);
and AND3 (N7042, N7032, N4420, N6168);
xor XOR2 (N7043, N7039, N4515);
nand NAND2 (N7044, N7023, N4667);
nor NOR4 (N7045, N7043, N4242, N801, N2029);
xor XOR2 (N7046, N7044, N2971);
nand NAND3 (N7047, N7034, N6350, N1351);
not NOT1 (N7048, N7041);
and AND4 (N7049, N7042, N2155, N6730, N180);
nand NAND4 (N7050, N7037, N3274, N2965, N5382);
nor NOR3 (N7051, N7047, N5433, N1621);
not NOT1 (N7052, N7031);
xor XOR2 (N7053, N7036, N3188);
buf BUF1 (N7054, N7045);
and AND2 (N7055, N7054, N6658);
not NOT1 (N7056, N7053);
and AND2 (N7057, N7048, N2188);
and AND3 (N7058, N7040, N901, N5687);
xor XOR2 (N7059, N7057, N5373);
nand NAND2 (N7060, N7055, N6259);
xor XOR2 (N7061, N7059, N2462);
nor NOR4 (N7062, N7038, N6671, N3169, N2914);
nor NOR4 (N7063, N7046, N6147, N1426, N6337);
nand NAND2 (N7064, N7061, N4822);
nand NAND4 (N7065, N7050, N2838, N2137, N535);
or OR2 (N7066, N7064, N2845);
xor XOR2 (N7067, N7058, N1397);
buf BUF1 (N7068, N7060);
buf BUF1 (N7069, N7052);
buf BUF1 (N7070, N7049);
and AND3 (N7071, N7068, N3252, N7005);
nor NOR3 (N7072, N7067, N3225, N1935);
nand NAND3 (N7073, N7051, N1184, N3395);
nand NAND3 (N7074, N7066, N532, N1607);
xor XOR2 (N7075, N7070, N6660);
not NOT1 (N7076, N7062);
nand NAND2 (N7077, N7065, N4798);
not NOT1 (N7078, N7072);
buf BUF1 (N7079, N7078);
and AND2 (N7080, N7076, N6905);
or OR4 (N7081, N7077, N5366, N432, N2812);
and AND4 (N7082, N7056, N4024, N1678, N1515);
buf BUF1 (N7083, N7075);
or OR4 (N7084, N7082, N3778, N1116, N2750);
and AND2 (N7085, N7063, N4570);
not NOT1 (N7086, N7073);
or OR2 (N7087, N7071, N2434);
xor XOR2 (N7088, N7080, N4023);
nor NOR3 (N7089, N7074, N6174, N6153);
nand NAND3 (N7090, N7088, N5273, N4712);
xor XOR2 (N7091, N7085, N7018);
not NOT1 (N7092, N7089);
xor XOR2 (N7093, N7091, N6604);
nand NAND4 (N7094, N7084, N6394, N6151, N2995);
nor NOR2 (N7095, N7093, N2896);
and AND2 (N7096, N7083, N2337);
or OR2 (N7097, N7079, N3444);
buf BUF1 (N7098, N7096);
nand NAND3 (N7099, N7090, N6227, N2713);
or OR4 (N7100, N7086, N6057, N4707, N1187);
nand NAND4 (N7101, N7095, N2788, N3256, N5003);
nand NAND3 (N7102, N7087, N458, N299);
and AND2 (N7103, N7102, N898);
not NOT1 (N7104, N7081);
not NOT1 (N7105, N7101);
buf BUF1 (N7106, N7105);
xor XOR2 (N7107, N7069, N4026);
nand NAND4 (N7108, N7098, N1124, N902, N5802);
nand NAND3 (N7109, N7094, N3667, N4467);
or OR4 (N7110, N7103, N3880, N4402, N1964);
not NOT1 (N7111, N7109);
buf BUF1 (N7112, N7106);
buf BUF1 (N7113, N7092);
xor XOR2 (N7114, N7099, N4456);
and AND3 (N7115, N7104, N5243, N4579);
and AND4 (N7116, N7100, N3244, N6729, N808);
xor XOR2 (N7117, N7115, N3113);
or OR2 (N7118, N7108, N6724);
and AND3 (N7119, N7118, N4509, N3184);
nor NOR2 (N7120, N7116, N923);
buf BUF1 (N7121, N7120);
nor NOR2 (N7122, N7114, N3063);
nand NAND4 (N7123, N7111, N5903, N4709, N2406);
and AND4 (N7124, N7121, N2395, N1931, N1162);
or OR2 (N7125, N7123, N6260);
not NOT1 (N7126, N7110);
or OR4 (N7127, N7097, N4903, N6435, N4960);
buf BUF1 (N7128, N7112);
nor NOR4 (N7129, N7119, N1468, N4304, N3347);
not NOT1 (N7130, N7117);
not NOT1 (N7131, N7126);
and AND2 (N7132, N7129, N1480);
and AND3 (N7133, N7125, N3128, N986);
xor XOR2 (N7134, N7127, N5401);
nand NAND3 (N7135, N7134, N754, N4308);
buf BUF1 (N7136, N7131);
nor NOR2 (N7137, N7128, N4646);
xor XOR2 (N7138, N7132, N4943);
or OR3 (N7139, N7122, N4860, N1699);
xor XOR2 (N7140, N7138, N2016);
and AND4 (N7141, N7140, N4878, N630, N7011);
or OR2 (N7142, N7135, N2019);
nand NAND4 (N7143, N7136, N1230, N3454, N1414);
nand NAND3 (N7144, N7137, N6833, N1021);
xor XOR2 (N7145, N7130, N512);
nand NAND2 (N7146, N7133, N1900);
or OR3 (N7147, N7142, N5311, N128);
not NOT1 (N7148, N7147);
not NOT1 (N7149, N7124);
and AND3 (N7150, N7146, N1621, N6749);
and AND4 (N7151, N7144, N252, N5824, N3657);
buf BUF1 (N7152, N7150);
not NOT1 (N7153, N7149);
not NOT1 (N7154, N7148);
nor NOR2 (N7155, N7153, N2415);
or OR3 (N7156, N7151, N3272, N4570);
or OR3 (N7157, N7139, N6116, N5510);
and AND2 (N7158, N7157, N1968);
not NOT1 (N7159, N7107);
not NOT1 (N7160, N7155);
and AND3 (N7161, N7154, N5225, N1665);
nand NAND4 (N7162, N7156, N2330, N2058, N7098);
nand NAND2 (N7163, N7113, N5974);
or OR2 (N7164, N7161, N3854);
xor XOR2 (N7165, N7164, N3377);
nor NOR4 (N7166, N7141, N4798, N1522, N3936);
and AND2 (N7167, N7158, N1242);
or OR4 (N7168, N7163, N4370, N4797, N4435);
not NOT1 (N7169, N7143);
buf BUF1 (N7170, N7162);
buf BUF1 (N7171, N7165);
or OR3 (N7172, N7170, N870, N4625);
or OR3 (N7173, N7145, N2932, N784);
or OR2 (N7174, N7168, N1290);
not NOT1 (N7175, N7172);
nand NAND4 (N7176, N7152, N5158, N3158, N469);
and AND2 (N7177, N7167, N5881);
xor XOR2 (N7178, N7175, N6958);
not NOT1 (N7179, N7171);
buf BUF1 (N7180, N7179);
xor XOR2 (N7181, N7180, N4285);
not NOT1 (N7182, N7173);
buf BUF1 (N7183, N7174);
xor XOR2 (N7184, N7182, N6418);
xor XOR2 (N7185, N7160, N2324);
and AND3 (N7186, N7183, N2690, N5642);
xor XOR2 (N7187, N7178, N1542);
nor NOR3 (N7188, N7159, N1022, N548);
nor NOR4 (N7189, N7181, N6487, N2508, N5804);
not NOT1 (N7190, N7189);
nand NAND3 (N7191, N7188, N3551, N6);
xor XOR2 (N7192, N7191, N5854);
nor NOR2 (N7193, N7176, N203);
nor NOR4 (N7194, N7185, N2323, N3920, N1720);
xor XOR2 (N7195, N7194, N1946);
and AND4 (N7196, N7193, N2506, N647, N561);
and AND3 (N7197, N7184, N4623, N5812);
or OR2 (N7198, N7166, N3918);
xor XOR2 (N7199, N7196, N863);
buf BUF1 (N7200, N7187);
nor NOR4 (N7201, N7195, N689, N3539, N1975);
not NOT1 (N7202, N7186);
nor NOR3 (N7203, N7201, N3084, N486);
nand NAND2 (N7204, N7200, N4505);
nor NOR3 (N7205, N7190, N6619, N1628);
xor XOR2 (N7206, N7202, N5085);
buf BUF1 (N7207, N7177);
nand NAND4 (N7208, N7169, N3209, N1863, N6829);
not NOT1 (N7209, N7205);
buf BUF1 (N7210, N7204);
buf BUF1 (N7211, N7208);
nand NAND4 (N7212, N7211, N2349, N6778, N6982);
xor XOR2 (N7213, N7198, N2523);
and AND3 (N7214, N7212, N3127, N320);
xor XOR2 (N7215, N7207, N937);
or OR3 (N7216, N7206, N4878, N3940);
xor XOR2 (N7217, N7214, N3208);
xor XOR2 (N7218, N7192, N1484);
not NOT1 (N7219, N7203);
or OR2 (N7220, N7210, N107);
or OR4 (N7221, N7218, N6495, N6150, N856);
nand NAND4 (N7222, N7199, N6458, N6620, N178);
nor NOR2 (N7223, N7197, N5441);
nor NOR3 (N7224, N7223, N3166, N4605);
or OR3 (N7225, N7220, N512, N3106);
buf BUF1 (N7226, N7217);
xor XOR2 (N7227, N7221, N4230);
and AND3 (N7228, N7227, N1877, N5308);
nor NOR3 (N7229, N7215, N2629, N2709);
xor XOR2 (N7230, N7224, N3774);
not NOT1 (N7231, N7228);
xor XOR2 (N7232, N7230, N1178);
nor NOR3 (N7233, N7229, N4587, N1913);
or OR4 (N7234, N7233, N5888, N2138, N1632);
nor NOR4 (N7235, N7209, N3875, N4309, N3323);
buf BUF1 (N7236, N7234);
not NOT1 (N7237, N7213);
nand NAND4 (N7238, N7222, N5501, N770, N306);
nand NAND3 (N7239, N7216, N2074, N6034);
nor NOR4 (N7240, N7238, N3281, N4263, N4294);
and AND3 (N7241, N7236, N4029, N5219);
nor NOR2 (N7242, N7239, N2886);
nand NAND2 (N7243, N7237, N3660);
or OR2 (N7244, N7240, N7236);
nor NOR3 (N7245, N7235, N3679, N1795);
nor NOR4 (N7246, N7232, N1056, N625, N1864);
or OR3 (N7247, N7246, N6210, N3886);
xor XOR2 (N7248, N7219, N1344);
not NOT1 (N7249, N7242);
nand NAND4 (N7250, N7247, N2971, N1826, N5112);
nor NOR2 (N7251, N7225, N864);
nand NAND4 (N7252, N7226, N6237, N6832, N448);
xor XOR2 (N7253, N7251, N2470);
nand NAND3 (N7254, N7248, N1366, N5469);
not NOT1 (N7255, N7244);
or OR2 (N7256, N7254, N494);
or OR3 (N7257, N7253, N5923, N6590);
buf BUF1 (N7258, N7257);
not NOT1 (N7259, N7245);
and AND4 (N7260, N7250, N2183, N3036, N1349);
or OR3 (N7261, N7241, N5218, N2373);
nor NOR2 (N7262, N7249, N648);
not NOT1 (N7263, N7259);
not NOT1 (N7264, N7262);
and AND2 (N7265, N7260, N2133);
or OR3 (N7266, N7256, N6470, N343);
buf BUF1 (N7267, N7252);
nor NOR3 (N7268, N7263, N6000, N3051);
nor NOR4 (N7269, N7267, N6113, N4457, N6347);
or OR2 (N7270, N7264, N254);
and AND3 (N7271, N7270, N5926, N5685);
nand NAND2 (N7272, N7231, N3323);
not NOT1 (N7273, N7272);
buf BUF1 (N7274, N7271);
xor XOR2 (N7275, N7269, N2060);
xor XOR2 (N7276, N7266, N909);
or OR4 (N7277, N7276, N1256, N2031, N3048);
nand NAND3 (N7278, N7277, N2257, N2519);
and AND2 (N7279, N7265, N4328);
nor NOR3 (N7280, N7255, N1666, N182);
or OR3 (N7281, N7280, N405, N4639);
xor XOR2 (N7282, N7261, N2853);
not NOT1 (N7283, N7282);
nand NAND2 (N7284, N7278, N6664);
nor NOR3 (N7285, N7283, N870, N5992);
not NOT1 (N7286, N7279);
buf BUF1 (N7287, N7281);
and AND4 (N7288, N7286, N4747, N3814, N5068);
not NOT1 (N7289, N7273);
buf BUF1 (N7290, N7287);
or OR3 (N7291, N7288, N1829, N4337);
xor XOR2 (N7292, N7290, N7106);
nor NOR2 (N7293, N7243, N1488);
nor NOR4 (N7294, N7293, N1651, N3455, N5443);
buf BUF1 (N7295, N7289);
nor NOR4 (N7296, N7285, N1878, N4580, N4726);
not NOT1 (N7297, N7274);
nand NAND4 (N7298, N7297, N6674, N4504, N7267);
nor NOR3 (N7299, N7292, N6007, N131);
or OR2 (N7300, N7284, N5956);
buf BUF1 (N7301, N7258);
buf BUF1 (N7302, N7299);
or OR2 (N7303, N7294, N5930);
or OR4 (N7304, N7268, N168, N3120, N2641);
buf BUF1 (N7305, N7301);
or OR3 (N7306, N7298, N2169, N3996);
and AND3 (N7307, N7295, N3687, N2906);
buf BUF1 (N7308, N7307);
nor NOR4 (N7309, N7308, N6601, N5432, N4663);
buf BUF1 (N7310, N7309);
nor NOR2 (N7311, N7300, N4521);
not NOT1 (N7312, N7310);
xor XOR2 (N7313, N7311, N6426);
or OR4 (N7314, N7302, N6874, N5384, N2077);
nor NOR3 (N7315, N7303, N5359, N7047);
nand NAND2 (N7316, N7312, N5758);
not NOT1 (N7317, N7305);
or OR2 (N7318, N7296, N3309);
and AND3 (N7319, N7291, N4266, N1208);
nand NAND4 (N7320, N7275, N6928, N3126, N4592);
and AND4 (N7321, N7319, N7304, N4634, N6881);
buf BUF1 (N7322, N4048);
not NOT1 (N7323, N7321);
not NOT1 (N7324, N7306);
nand NAND3 (N7325, N7323, N2021, N5146);
buf BUF1 (N7326, N7313);
buf BUF1 (N7327, N7326);
not NOT1 (N7328, N7316);
buf BUF1 (N7329, N7328);
buf BUF1 (N7330, N7324);
and AND3 (N7331, N7322, N428, N3624);
nand NAND2 (N7332, N7315, N2015);
not NOT1 (N7333, N7320);
nor NOR2 (N7334, N7329, N253);
xor XOR2 (N7335, N7314, N2492);
xor XOR2 (N7336, N7330, N2992);
or OR3 (N7337, N7317, N7197, N5362);
and AND4 (N7338, N7318, N7100, N2724, N3007);
nor NOR2 (N7339, N7331, N1173);
nor NOR4 (N7340, N7337, N3184, N6504, N7175);
or OR2 (N7341, N7336, N1608);
buf BUF1 (N7342, N7327);
and AND2 (N7343, N7341, N4710);
xor XOR2 (N7344, N7340, N201);
nor NOR4 (N7345, N7339, N6570, N7342, N4758);
buf BUF1 (N7346, N3586);
or OR3 (N7347, N7345, N415, N3348);
or OR3 (N7348, N7346, N6353, N2789);
or OR4 (N7349, N7347, N939, N4971, N2148);
or OR4 (N7350, N7325, N1875, N1102, N4671);
or OR2 (N7351, N7349, N1898);
not NOT1 (N7352, N7351);
xor XOR2 (N7353, N7348, N1032);
or OR4 (N7354, N7343, N1040, N4261, N4304);
buf BUF1 (N7355, N7344);
nor NOR4 (N7356, N7352, N4729, N2661, N5862);
nand NAND2 (N7357, N7355, N1464);
buf BUF1 (N7358, N7332);
or OR4 (N7359, N7338, N4168, N4771, N1485);
nor NOR3 (N7360, N7334, N5590, N2127);
nor NOR3 (N7361, N7360, N1918, N6893);
and AND4 (N7362, N7359, N2019, N2410, N3650);
not NOT1 (N7363, N7357);
and AND3 (N7364, N7358, N5452, N5256);
nand NAND3 (N7365, N7353, N743, N5590);
or OR2 (N7366, N7365, N1286);
buf BUF1 (N7367, N7335);
or OR3 (N7368, N7361, N3618, N3150);
nor NOR2 (N7369, N7333, N6128);
buf BUF1 (N7370, N7362);
not NOT1 (N7371, N7367);
buf BUF1 (N7372, N7371);
xor XOR2 (N7373, N7370, N3773);
buf BUF1 (N7374, N7363);
and AND2 (N7375, N7372, N2031);
nand NAND4 (N7376, N7374, N4613, N5726, N1322);
and AND4 (N7377, N7350, N5214, N7295, N2736);
nor NOR3 (N7378, N7369, N2988, N2369);
xor XOR2 (N7379, N7377, N4897);
xor XOR2 (N7380, N7364, N461);
buf BUF1 (N7381, N7379);
nand NAND2 (N7382, N7375, N994);
or OR3 (N7383, N7382, N1670, N2583);
nor NOR2 (N7384, N7383, N1748);
nand NAND2 (N7385, N7366, N857);
not NOT1 (N7386, N7385);
xor XOR2 (N7387, N7373, N4575);
buf BUF1 (N7388, N7384);
xor XOR2 (N7389, N7386, N7046);
nor NOR3 (N7390, N7354, N1450, N5311);
and AND3 (N7391, N7388, N3956, N3932);
xor XOR2 (N7392, N7356, N6926);
not NOT1 (N7393, N7389);
or OR2 (N7394, N7376, N154);
buf BUF1 (N7395, N7390);
nand NAND3 (N7396, N7368, N6073, N1225);
nand NAND4 (N7397, N7396, N2584, N6167, N2041);
or OR4 (N7398, N7392, N6083, N2472, N5445);
and AND3 (N7399, N7391, N4710, N1360);
nor NOR3 (N7400, N7380, N3805, N2688);
xor XOR2 (N7401, N7378, N5646);
buf BUF1 (N7402, N7395);
xor XOR2 (N7403, N7400, N3046);
nand NAND2 (N7404, N7401, N2136);
or OR3 (N7405, N7402, N3720, N5337);
not NOT1 (N7406, N7404);
not NOT1 (N7407, N7397);
or OR2 (N7408, N7403, N325);
buf BUF1 (N7409, N7407);
nor NOR2 (N7410, N7405, N1596);
nand NAND2 (N7411, N7398, N5622);
or OR4 (N7412, N7411, N3263, N1603, N3342);
xor XOR2 (N7413, N7408, N7226);
buf BUF1 (N7414, N7393);
nand NAND4 (N7415, N7387, N5973, N6626, N4740);
nor NOR4 (N7416, N7394, N7338, N7088, N4370);
or OR4 (N7417, N7406, N3679, N6418, N5731);
and AND4 (N7418, N7413, N1147, N5525, N1549);
or OR3 (N7419, N7412, N6886, N5918);
and AND3 (N7420, N7399, N7122, N4500);
xor XOR2 (N7421, N7410, N7340);
not NOT1 (N7422, N7414);
xor XOR2 (N7423, N7418, N3210);
and AND2 (N7424, N7415, N1119);
buf BUF1 (N7425, N7422);
not NOT1 (N7426, N7425);
buf BUF1 (N7427, N7420);
buf BUF1 (N7428, N7424);
not NOT1 (N7429, N7417);
or OR3 (N7430, N7429, N1304, N5010);
nor NOR2 (N7431, N7426, N3712);
xor XOR2 (N7432, N7381, N7259);
and AND3 (N7433, N7421, N3886, N1846);
not NOT1 (N7434, N7409);
or OR2 (N7435, N7427, N3516);
or OR4 (N7436, N7435, N5841, N7071, N3599);
and AND4 (N7437, N7423, N949, N3968, N3924);
nor NOR3 (N7438, N7434, N1490, N4073);
not NOT1 (N7439, N7432);
or OR4 (N7440, N7436, N6295, N5066, N5818);
or OR4 (N7441, N7439, N979, N6342, N798);
or OR2 (N7442, N7430, N5474);
buf BUF1 (N7443, N7433);
not NOT1 (N7444, N7438);
nor NOR4 (N7445, N7441, N4579, N6795, N4743);
or OR4 (N7446, N7444, N3568, N624, N2162);
or OR4 (N7447, N7445, N1590, N1375, N5197);
xor XOR2 (N7448, N7437, N5081);
nand NAND3 (N7449, N7447, N5797, N5690);
and AND2 (N7450, N7443, N1495);
xor XOR2 (N7451, N7428, N1042);
or OR4 (N7452, N7450, N4177, N3828, N3275);
not NOT1 (N7453, N7451);
nor NOR3 (N7454, N7452, N3648, N803);
nor NOR4 (N7455, N7440, N2362, N2959, N1066);
nor NOR4 (N7456, N7453, N5177, N3752, N5587);
nand NAND3 (N7457, N7454, N2148, N5355);
and AND4 (N7458, N7449, N4496, N4148, N1685);
and AND3 (N7459, N7431, N2255, N2803);
nand NAND4 (N7460, N7458, N7189, N2851, N6522);
or OR3 (N7461, N7448, N4192, N2249);
and AND4 (N7462, N7419, N1748, N5294, N3516);
or OR2 (N7463, N7442, N966);
or OR3 (N7464, N7416, N6476, N4737);
xor XOR2 (N7465, N7463, N6990);
and AND3 (N7466, N7461, N5314, N1497);
nand NAND2 (N7467, N7459, N4768);
buf BUF1 (N7468, N7467);
or OR3 (N7469, N7460, N6392, N437);
and AND2 (N7470, N7465, N6825);
and AND2 (N7471, N7464, N7305);
and AND4 (N7472, N7462, N4758, N501, N7055);
xor XOR2 (N7473, N7457, N6852);
or OR2 (N7474, N7470, N4400);
buf BUF1 (N7475, N7473);
nor NOR4 (N7476, N7468, N5712, N5690, N4618);
not NOT1 (N7477, N7471);
and AND2 (N7478, N7469, N7221);
buf BUF1 (N7479, N7474);
and AND2 (N7480, N7475, N5327);
nor NOR4 (N7481, N7477, N5267, N854, N45);
nand NAND4 (N7482, N7456, N3750, N2798, N2111);
and AND3 (N7483, N7480, N612, N5956);
nand NAND3 (N7484, N7446, N1884, N7346);
nand NAND4 (N7485, N7479, N1029, N1026, N5021);
or OR4 (N7486, N7484, N3713, N1834, N3864);
or OR3 (N7487, N7466, N6323, N1744);
or OR3 (N7488, N7485, N7013, N2055);
or OR4 (N7489, N7483, N1284, N1576, N1548);
nor NOR2 (N7490, N7481, N5674);
buf BUF1 (N7491, N7490);
not NOT1 (N7492, N7455);
buf BUF1 (N7493, N7492);
and AND4 (N7494, N7476, N5403, N2282, N6340);
and AND4 (N7495, N7486, N1077, N5292, N6523);
and AND4 (N7496, N7478, N4081, N4884, N6143);
not NOT1 (N7497, N7496);
xor XOR2 (N7498, N7482, N6192);
not NOT1 (N7499, N7488);
nor NOR4 (N7500, N7487, N4933, N6990, N6564);
nand NAND2 (N7501, N7495, N5519);
nand NAND3 (N7502, N7497, N2307, N7273);
not NOT1 (N7503, N7502);
nor NOR3 (N7504, N7472, N4773, N2152);
xor XOR2 (N7505, N7504, N1660);
and AND2 (N7506, N7500, N6274);
and AND4 (N7507, N7506, N3056, N5598, N979);
nor NOR3 (N7508, N7498, N6256, N2329);
nor NOR3 (N7509, N7508, N4377, N2789);
xor XOR2 (N7510, N7503, N5600);
or OR2 (N7511, N7493, N1742);
or OR4 (N7512, N7499, N4658, N5411, N2127);
buf BUF1 (N7513, N7509);
nand NAND4 (N7514, N7501, N3416, N5938, N5071);
nand NAND3 (N7515, N7494, N190, N1492);
nor NOR4 (N7516, N7510, N2677, N3929, N5583);
nor NOR3 (N7517, N7489, N2962, N3974);
and AND2 (N7518, N7491, N5347);
not NOT1 (N7519, N7518);
buf BUF1 (N7520, N7519);
nand NAND2 (N7521, N7512, N5254);
nor NOR3 (N7522, N7520, N4439, N1038);
nand NAND4 (N7523, N7516, N331, N4267, N588);
buf BUF1 (N7524, N7505);
xor XOR2 (N7525, N7524, N5671);
or OR4 (N7526, N7517, N4047, N7240, N5151);
or OR3 (N7527, N7514, N6107, N4205);
nor NOR3 (N7528, N7515, N1372, N773);
xor XOR2 (N7529, N7526, N1085);
and AND4 (N7530, N7527, N298, N4740, N4380);
or OR2 (N7531, N7529, N2090);
xor XOR2 (N7532, N7511, N6538);
nor NOR3 (N7533, N7513, N5905, N6987);
or OR2 (N7534, N7525, N6089);
nand NAND3 (N7535, N7530, N1575, N685);
not NOT1 (N7536, N7521);
nand NAND2 (N7537, N7507, N2143);
nor NOR3 (N7538, N7523, N4822, N1204);
buf BUF1 (N7539, N7535);
buf BUF1 (N7540, N7536);
nand NAND4 (N7541, N7538, N3242, N3064, N274);
nand NAND2 (N7542, N7541, N1120);
and AND3 (N7543, N7528, N803, N3312);
not NOT1 (N7544, N7540);
buf BUF1 (N7545, N7544);
buf BUF1 (N7546, N7533);
nor NOR2 (N7547, N7534, N6749);
and AND2 (N7548, N7547, N1544);
buf BUF1 (N7549, N7539);
buf BUF1 (N7550, N7542);
xor XOR2 (N7551, N7522, N6961);
nand NAND2 (N7552, N7532, N2405);
buf BUF1 (N7553, N7550);
not NOT1 (N7554, N7548);
buf BUF1 (N7555, N7537);
buf BUF1 (N7556, N7549);
buf BUF1 (N7557, N7556);
xor XOR2 (N7558, N7554, N5184);
buf BUF1 (N7559, N7558);
buf BUF1 (N7560, N7553);
or OR4 (N7561, N7552, N1864, N6979, N2880);
not NOT1 (N7562, N7561);
nor NOR3 (N7563, N7543, N186, N3807);
nand NAND4 (N7564, N7559, N7000, N5784, N7193);
not NOT1 (N7565, N7555);
not NOT1 (N7566, N7563);
buf BUF1 (N7567, N7546);
not NOT1 (N7568, N7566);
buf BUF1 (N7569, N7564);
nor NOR4 (N7570, N7560, N2537, N7348, N6753);
buf BUF1 (N7571, N7551);
and AND4 (N7572, N7570, N718, N3012, N3581);
and AND2 (N7573, N7531, N7504);
and AND3 (N7574, N7572, N6446, N685);
buf BUF1 (N7575, N7569);
and AND4 (N7576, N7562, N4180, N2810, N3068);
and AND2 (N7577, N7568, N4103);
and AND2 (N7578, N7577, N2667);
not NOT1 (N7579, N7571);
buf BUF1 (N7580, N7565);
or OR4 (N7581, N7574, N5100, N5525, N2495);
and AND4 (N7582, N7579, N5009, N5594, N4894);
nor NOR4 (N7583, N7545, N7375, N6592, N6886);
not NOT1 (N7584, N7581);
and AND2 (N7585, N7582, N193);
nand NAND2 (N7586, N7585, N4999);
nand NAND4 (N7587, N7586, N4994, N2386, N6948);
nand NAND4 (N7588, N7573, N867, N6491, N6696);
xor XOR2 (N7589, N7575, N4142);
or OR3 (N7590, N7583, N516, N3063);
not NOT1 (N7591, N7587);
buf BUF1 (N7592, N7580);
and AND2 (N7593, N7589, N6669);
and AND4 (N7594, N7590, N7492, N1294, N5394);
not NOT1 (N7595, N7591);
nor NOR2 (N7596, N7594, N4819);
nand NAND2 (N7597, N7588, N748);
or OR3 (N7598, N7592, N6613, N2850);
xor XOR2 (N7599, N7584, N3477);
xor XOR2 (N7600, N7593, N3366);
xor XOR2 (N7601, N7596, N136);
and AND4 (N7602, N7601, N6333, N7081, N3273);
nor NOR3 (N7603, N7595, N5239, N1578);
or OR3 (N7604, N7576, N1286, N3593);
xor XOR2 (N7605, N7603, N3118);
not NOT1 (N7606, N7604);
or OR2 (N7607, N7598, N5603);
nor NOR3 (N7608, N7599, N7355, N1873);
not NOT1 (N7609, N7578);
nor NOR2 (N7610, N7600, N6994);
xor XOR2 (N7611, N7602, N6226);
not NOT1 (N7612, N7609);
and AND3 (N7613, N7605, N7545, N3880);
not NOT1 (N7614, N7612);
and AND4 (N7615, N7557, N5990, N868, N6875);
not NOT1 (N7616, N7614);
buf BUF1 (N7617, N7613);
nor NOR2 (N7618, N7610, N820);
buf BUF1 (N7619, N7606);
nor NOR4 (N7620, N7608, N2986, N449, N1808);
buf BUF1 (N7621, N7617);
xor XOR2 (N7622, N7567, N4499);
xor XOR2 (N7623, N7618, N6534);
and AND4 (N7624, N7622, N5870, N1630, N7434);
nor NOR2 (N7625, N7621, N5036);
nor NOR4 (N7626, N7619, N7020, N4267, N32);
nor NOR4 (N7627, N7624, N7057, N4917, N2998);
nor NOR4 (N7628, N7616, N5348, N1152, N2879);
nand NAND4 (N7629, N7611, N3949, N3970, N474);
xor XOR2 (N7630, N7607, N6690);
nor NOR4 (N7631, N7627, N3776, N6330, N4364);
buf BUF1 (N7632, N7628);
buf BUF1 (N7633, N7629);
nor NOR4 (N7634, N7623, N5135, N6517, N1389);
nand NAND3 (N7635, N7634, N7035, N6895);
or OR4 (N7636, N7631, N881, N795, N7320);
nand NAND3 (N7637, N7597, N593, N4946);
or OR3 (N7638, N7615, N1126, N4707);
or OR3 (N7639, N7637, N7307, N1143);
not NOT1 (N7640, N7636);
buf BUF1 (N7641, N7638);
or OR3 (N7642, N7625, N360, N6461);
not NOT1 (N7643, N7620);
xor XOR2 (N7644, N7643, N4793);
or OR2 (N7645, N7626, N511);
not NOT1 (N7646, N7639);
or OR4 (N7647, N7633, N6461, N3456, N7434);
and AND2 (N7648, N7645, N5745);
buf BUF1 (N7649, N7647);
or OR3 (N7650, N7630, N6313, N4503);
nor NOR3 (N7651, N7641, N2209, N2961);
and AND3 (N7652, N7649, N196, N6710);
xor XOR2 (N7653, N7652, N700);
or OR4 (N7654, N7640, N3639, N5703, N3172);
nor NOR2 (N7655, N7632, N1312);
xor XOR2 (N7656, N7654, N6942);
buf BUF1 (N7657, N7656);
nand NAND3 (N7658, N7655, N1023, N5645);
and AND2 (N7659, N7653, N6427);
xor XOR2 (N7660, N7648, N7332);
or OR3 (N7661, N7651, N3933, N7595);
or OR3 (N7662, N7646, N3527, N6599);
nor NOR4 (N7663, N7642, N2391, N112, N7657);
nor NOR4 (N7664, N1838, N2769, N5131, N1392);
not NOT1 (N7665, N7635);
not NOT1 (N7666, N7663);
and AND2 (N7667, N7666, N5200);
xor XOR2 (N7668, N7660, N3632);
buf BUF1 (N7669, N7665);
or OR3 (N7670, N7659, N7089, N1771);
buf BUF1 (N7671, N7667);
and AND2 (N7672, N7650, N1851);
nor NOR3 (N7673, N7662, N2896, N975);
and AND2 (N7674, N7673, N2844);
nand NAND2 (N7675, N7669, N4610);
nand NAND4 (N7676, N7664, N286, N501, N101);
xor XOR2 (N7677, N7670, N5359);
or OR3 (N7678, N7674, N1941, N784);
not NOT1 (N7679, N7676);
nor NOR2 (N7680, N7668, N1030);
or OR2 (N7681, N7675, N3051);
not NOT1 (N7682, N7681);
nor NOR3 (N7683, N7682, N2352, N5481);
and AND3 (N7684, N7658, N648, N7576);
buf BUF1 (N7685, N7679);
xor XOR2 (N7686, N7680, N3418);
nand NAND2 (N7687, N7661, N3115);
xor XOR2 (N7688, N7684, N759);
not NOT1 (N7689, N7671);
and AND2 (N7690, N7677, N4640);
nand NAND4 (N7691, N7672, N6018, N915, N2610);
nor NOR3 (N7692, N7691, N3797, N1196);
not NOT1 (N7693, N7688);
buf BUF1 (N7694, N7687);
or OR4 (N7695, N7694, N416, N5639, N5243);
not NOT1 (N7696, N7695);
nor NOR3 (N7697, N7689, N4015, N6386);
nand NAND3 (N7698, N7697, N3737, N172);
xor XOR2 (N7699, N7696, N2584);
or OR4 (N7700, N7685, N951, N2251, N6853);
buf BUF1 (N7701, N7690);
not NOT1 (N7702, N7683);
and AND4 (N7703, N7702, N1606, N855, N5469);
buf BUF1 (N7704, N7686);
or OR4 (N7705, N7692, N997, N1177, N3331);
xor XOR2 (N7706, N7704, N5901);
nor NOR3 (N7707, N7700, N6706, N5803);
and AND2 (N7708, N7703, N1438);
xor XOR2 (N7709, N7678, N4429);
nor NOR4 (N7710, N7701, N120, N2294, N3945);
and AND2 (N7711, N7698, N5737);
and AND4 (N7712, N7709, N5311, N1118, N729);
or OR3 (N7713, N7706, N4144, N3416);
or OR2 (N7714, N7707, N1357);
not NOT1 (N7715, N7705);
xor XOR2 (N7716, N7713, N6301);
buf BUF1 (N7717, N7712);
buf BUF1 (N7718, N7710);
nand NAND3 (N7719, N7717, N2551, N3351);
buf BUF1 (N7720, N7715);
buf BUF1 (N7721, N7714);
buf BUF1 (N7722, N7718);
and AND2 (N7723, N7644, N3815);
nand NAND2 (N7724, N7722, N4369);
nor NOR3 (N7725, N7719, N4144, N7603);
or OR3 (N7726, N7720, N6146, N1539);
and AND4 (N7727, N7699, N6882, N2627, N4011);
not NOT1 (N7728, N7724);
and AND2 (N7729, N7726, N3715);
or OR4 (N7730, N7721, N137, N818, N4555);
xor XOR2 (N7731, N7711, N4933);
xor XOR2 (N7732, N7730, N5629);
buf BUF1 (N7733, N7716);
or OR2 (N7734, N7729, N6442);
nand NAND2 (N7735, N7725, N4348);
nand NAND2 (N7736, N7734, N2240);
or OR2 (N7737, N7736, N6303);
buf BUF1 (N7738, N7727);
buf BUF1 (N7739, N7708);
and AND4 (N7740, N7739, N6218, N714, N5917);
xor XOR2 (N7741, N7738, N7237);
not NOT1 (N7742, N7733);
buf BUF1 (N7743, N7740);
nor NOR3 (N7744, N7742, N6153, N4334);
or OR3 (N7745, N7732, N1351, N1299);
and AND4 (N7746, N7723, N3575, N1007, N3648);
buf BUF1 (N7747, N7728);
nor NOR3 (N7748, N7735, N7745, N7588);
and AND4 (N7749, N2461, N6182, N3400, N699);
nor NOR3 (N7750, N7749, N1880, N7093);
and AND4 (N7751, N7693, N407, N219, N6131);
nand NAND3 (N7752, N7741, N788, N7133);
buf BUF1 (N7753, N7747);
buf BUF1 (N7754, N7751);
nand NAND4 (N7755, N7731, N6761, N6732, N2081);
or OR2 (N7756, N7753, N2389);
not NOT1 (N7757, N7748);
nor NOR4 (N7758, N7750, N4226, N3061, N3969);
not NOT1 (N7759, N7752);
or OR3 (N7760, N7757, N5109, N7674);
buf BUF1 (N7761, N7759);
nor NOR3 (N7762, N7737, N2430, N3839);
buf BUF1 (N7763, N7758);
not NOT1 (N7764, N7760);
and AND3 (N7765, N7764, N3502, N4593);
nor NOR3 (N7766, N7756, N6261, N2806);
xor XOR2 (N7767, N7746, N7736);
nor NOR2 (N7768, N7754, N7055);
or OR3 (N7769, N7766, N1047, N665);
nand NAND3 (N7770, N7761, N1089, N4761);
xor XOR2 (N7771, N7765, N4188);
nand NAND2 (N7772, N7743, N3175);
nor NOR2 (N7773, N7744, N7145);
and AND3 (N7774, N7769, N1072, N4618);
xor XOR2 (N7775, N7762, N7764);
nor NOR3 (N7776, N7774, N4860, N5236);
and AND4 (N7777, N7768, N3715, N529, N1738);
nor NOR2 (N7778, N7755, N7334);
and AND2 (N7779, N7777, N7142);
or OR4 (N7780, N7770, N6805, N5131, N2998);
nor NOR2 (N7781, N7767, N7488);
and AND2 (N7782, N7779, N3712);
nand NAND3 (N7783, N7771, N7525, N636);
not NOT1 (N7784, N7775);
or OR2 (N7785, N7780, N6099);
nor NOR4 (N7786, N7783, N6778, N5633, N1552);
nor NOR3 (N7787, N7776, N7178, N4370);
buf BUF1 (N7788, N7763);
nand NAND3 (N7789, N7778, N1868, N793);
or OR4 (N7790, N7788, N457, N137, N2492);
and AND3 (N7791, N7782, N5650, N1095);
nand NAND3 (N7792, N7791, N3544, N1345);
nand NAND4 (N7793, N7785, N118, N4605, N3142);
and AND3 (N7794, N7787, N3613, N1826);
not NOT1 (N7795, N7790);
nor NOR3 (N7796, N7789, N5451, N7334);
or OR4 (N7797, N7792, N3127, N5310, N4670);
and AND4 (N7798, N7794, N3417, N2749, N2769);
not NOT1 (N7799, N7786);
or OR3 (N7800, N7799, N2058, N1157);
not NOT1 (N7801, N7797);
and AND2 (N7802, N7798, N2858);
or OR3 (N7803, N7793, N956, N4206);
buf BUF1 (N7804, N7800);
and AND4 (N7805, N7803, N5101, N2546, N231);
or OR3 (N7806, N7801, N5611, N5006);
xor XOR2 (N7807, N7795, N5183);
and AND3 (N7808, N7784, N4972, N2989);
not NOT1 (N7809, N7804);
buf BUF1 (N7810, N7807);
xor XOR2 (N7811, N7796, N5221);
or OR4 (N7812, N7811, N217, N128, N6568);
or OR4 (N7813, N7812, N6233, N1649, N7559);
buf BUF1 (N7814, N7808);
nand NAND2 (N7815, N7781, N5052);
and AND3 (N7816, N7813, N5323, N5723);
nor NOR2 (N7817, N7814, N1295);
and AND3 (N7818, N7815, N4137, N7651);
buf BUF1 (N7819, N7805);
nor NOR4 (N7820, N7809, N5352, N2818, N2386);
nor NOR2 (N7821, N7816, N6676);
or OR3 (N7822, N7817, N7393, N6324);
nor NOR2 (N7823, N7818, N7028);
nand NAND2 (N7824, N7772, N1085);
xor XOR2 (N7825, N7820, N316);
or OR2 (N7826, N7821, N2182);
or OR3 (N7827, N7822, N7519, N2959);
and AND2 (N7828, N7819, N2863);
xor XOR2 (N7829, N7825, N5320);
nand NAND2 (N7830, N7826, N5412);
and AND2 (N7831, N7823, N238);
and AND3 (N7832, N7827, N2594, N1705);
nor NOR2 (N7833, N7828, N6484);
nand NAND4 (N7834, N7831, N6619, N7042, N956);
xor XOR2 (N7835, N7810, N4212);
not NOT1 (N7836, N7829);
nor NOR3 (N7837, N7832, N7423, N4457);
not NOT1 (N7838, N7773);
xor XOR2 (N7839, N7802, N6600);
or OR2 (N7840, N7836, N496);
not NOT1 (N7841, N7838);
nor NOR2 (N7842, N7834, N4799);
nor NOR4 (N7843, N7806, N3159, N2856, N4676);
not NOT1 (N7844, N7842);
nand NAND3 (N7845, N7840, N1357, N2000);
xor XOR2 (N7846, N7839, N1154);
and AND4 (N7847, N7824, N1569, N1631, N3069);
or OR2 (N7848, N7846, N7529);
buf BUF1 (N7849, N7833);
xor XOR2 (N7850, N7849, N4593);
and AND4 (N7851, N7845, N983, N5451, N4288);
nor NOR2 (N7852, N7841, N777);
or OR3 (N7853, N7851, N6114, N4600);
buf BUF1 (N7854, N7848);
xor XOR2 (N7855, N7835, N2173);
or OR2 (N7856, N7850, N7631);
nor NOR3 (N7857, N7853, N3587, N6292);
nor NOR2 (N7858, N7857, N4284);
nand NAND4 (N7859, N7844, N6566, N2978, N4918);
buf BUF1 (N7860, N7852);
or OR2 (N7861, N7860, N2375);
and AND4 (N7862, N7858, N3963, N1409, N5016);
xor XOR2 (N7863, N7861, N2827);
nor NOR2 (N7864, N7856, N1417);
and AND4 (N7865, N7847, N5979, N1141, N4275);
or OR2 (N7866, N7855, N5206);
nor NOR2 (N7867, N7864, N7719);
or OR3 (N7868, N7837, N5375, N7725);
xor XOR2 (N7869, N7862, N2873);
not NOT1 (N7870, N7867);
and AND4 (N7871, N7843, N1326, N4026, N3758);
and AND2 (N7872, N7868, N7835);
nor NOR3 (N7873, N7830, N5143, N49);
or OR4 (N7874, N7865, N6448, N2838, N1737);
nor NOR2 (N7875, N7859, N631);
xor XOR2 (N7876, N7863, N5972);
and AND3 (N7877, N7873, N3040, N6518);
nor NOR4 (N7878, N7876, N2687, N4474, N3665);
nor NOR2 (N7879, N7870, N6697);
and AND3 (N7880, N7875, N6124, N2526);
nand NAND2 (N7881, N7871, N2970);
or OR2 (N7882, N7866, N6089);
and AND4 (N7883, N7874, N5947, N7410, N5605);
nand NAND3 (N7884, N7880, N4956, N70);
or OR4 (N7885, N7854, N585, N4031, N758);
and AND4 (N7886, N7869, N7069, N1752, N4021);
nand NAND3 (N7887, N7886, N5237, N1296);
not NOT1 (N7888, N7872);
not NOT1 (N7889, N7887);
xor XOR2 (N7890, N7889, N7484);
or OR2 (N7891, N7883, N5671);
and AND3 (N7892, N7888, N7529, N998);
buf BUF1 (N7893, N7885);
buf BUF1 (N7894, N7878);
nand NAND2 (N7895, N7882, N4682);
xor XOR2 (N7896, N7877, N5506);
nand NAND3 (N7897, N7884, N6570, N3668);
nand NAND2 (N7898, N7896, N6875);
xor XOR2 (N7899, N7893, N6024);
or OR3 (N7900, N7894, N5591, N5457);
xor XOR2 (N7901, N7890, N3087);
xor XOR2 (N7902, N7891, N2991);
nand NAND2 (N7903, N7881, N6788);
not NOT1 (N7904, N7897);
not NOT1 (N7905, N7899);
nand NAND2 (N7906, N7902, N4105);
and AND4 (N7907, N7903, N1484, N2070, N4339);
or OR3 (N7908, N7905, N1656, N1172);
not NOT1 (N7909, N7901);
and AND2 (N7910, N7898, N1537);
xor XOR2 (N7911, N7879, N7489);
not NOT1 (N7912, N7904);
buf BUF1 (N7913, N7895);
not NOT1 (N7914, N7906);
not NOT1 (N7915, N7910);
nand NAND3 (N7916, N7909, N4176, N2855);
nand NAND2 (N7917, N7912, N4002);
buf BUF1 (N7918, N7900);
and AND3 (N7919, N7918, N3356, N7901);
nand NAND2 (N7920, N7917, N5287);
and AND4 (N7921, N7911, N1275, N1797, N230);
not NOT1 (N7922, N7920);
xor XOR2 (N7923, N7892, N2909);
nand NAND2 (N7924, N7914, N2916);
not NOT1 (N7925, N7921);
or OR3 (N7926, N7919, N6582, N7193);
nor NOR2 (N7927, N7913, N1239);
buf BUF1 (N7928, N7927);
not NOT1 (N7929, N7908);
xor XOR2 (N7930, N7922, N6797);
nor NOR2 (N7931, N7923, N64);
nand NAND4 (N7932, N7928, N1475, N778, N3999);
nand NAND3 (N7933, N7915, N340, N5004);
and AND4 (N7934, N7925, N5022, N1317, N2824);
xor XOR2 (N7935, N7926, N884);
nand NAND3 (N7936, N7933, N6229, N3765);
xor XOR2 (N7937, N7936, N4673);
buf BUF1 (N7938, N7935);
nand NAND3 (N7939, N7929, N5163, N7872);
not NOT1 (N7940, N7930);
nor NOR3 (N7941, N7934, N2764, N7437);
and AND4 (N7942, N7932, N3024, N236, N5460);
nor NOR3 (N7943, N7940, N5496, N3516);
xor XOR2 (N7944, N7924, N7288);
not NOT1 (N7945, N7941);
not NOT1 (N7946, N7943);
buf BUF1 (N7947, N7939);
buf BUF1 (N7948, N7945);
not NOT1 (N7949, N7942);
xor XOR2 (N7950, N7931, N1756);
nor NOR3 (N7951, N7916, N6653, N6447);
and AND3 (N7952, N7949, N643, N6851);
not NOT1 (N7953, N7952);
and AND3 (N7954, N7948, N5426, N3372);
and AND2 (N7955, N7950, N1055);
buf BUF1 (N7956, N7938);
nor NOR3 (N7957, N7954, N3506, N1859);
nor NOR2 (N7958, N7946, N93);
xor XOR2 (N7959, N7937, N3632);
not NOT1 (N7960, N7956);
not NOT1 (N7961, N7955);
xor XOR2 (N7962, N7944, N1816);
xor XOR2 (N7963, N7960, N1766);
buf BUF1 (N7964, N7958);
nor NOR2 (N7965, N7947, N4015);
or OR4 (N7966, N7961, N7210, N4045, N5612);
buf BUF1 (N7967, N7962);
and AND3 (N7968, N7966, N2645, N5397);
nand NAND3 (N7969, N7957, N7143, N6464);
nand NAND3 (N7970, N7907, N6687, N2870);
buf BUF1 (N7971, N7959);
nand NAND3 (N7972, N7969, N7600, N1241);
xor XOR2 (N7973, N7970, N30);
xor XOR2 (N7974, N7971, N3730);
xor XOR2 (N7975, N7951, N5198);
buf BUF1 (N7976, N7964);
nand NAND3 (N7977, N7973, N2804, N3451);
or OR4 (N7978, N7967, N6825, N3676, N6036);
and AND2 (N7979, N7974, N561);
nand NAND2 (N7980, N7975, N2193);
nand NAND4 (N7981, N7976, N542, N4627, N2395);
xor XOR2 (N7982, N7972, N2591);
nand NAND3 (N7983, N7978, N7370, N1464);
nor NOR2 (N7984, N7981, N4245);
not NOT1 (N7985, N7977);
nand NAND4 (N7986, N7968, N2268, N6602, N1357);
and AND2 (N7987, N7983, N4803);
or OR3 (N7988, N7984, N3710, N81);
buf BUF1 (N7989, N7982);
nand NAND3 (N7990, N7979, N7112, N7802);
xor XOR2 (N7991, N7987, N2340);
not NOT1 (N7992, N7965);
or OR2 (N7993, N7989, N841);
and AND4 (N7994, N7991, N1497, N1043, N4425);
not NOT1 (N7995, N7992);
xor XOR2 (N7996, N7986, N1941);
not NOT1 (N7997, N7985);
nand NAND4 (N7998, N7995, N3659, N4102, N5515);
and AND4 (N7999, N7994, N232, N7823, N2640);
nor NOR2 (N8000, N7990, N7996);
xor XOR2 (N8001, N7722, N2922);
nand NAND2 (N8002, N7988, N1225);
buf BUF1 (N8003, N8000);
xor XOR2 (N8004, N7999, N7248);
xor XOR2 (N8005, N8002, N3376);
not NOT1 (N8006, N7997);
xor XOR2 (N8007, N7953, N5354);
nor NOR4 (N8008, N8001, N4351, N7328, N5936);
nor NOR3 (N8009, N7963, N5422, N1287);
nand NAND4 (N8010, N8009, N1683, N483, N3794);
nor NOR3 (N8011, N8003, N3386, N459);
or OR4 (N8012, N8008, N371, N6731, N7262);
and AND3 (N8013, N7980, N261, N5816);
nand NAND2 (N8014, N8011, N6597);
and AND2 (N8015, N8014, N6372);
or OR3 (N8016, N8013, N1541, N7088);
not NOT1 (N8017, N8004);
buf BUF1 (N8018, N8007);
endmodule