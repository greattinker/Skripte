// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17;

output N914,N913,N910,N897,N915,N888,N916,N900,N903,N917;

or OR3 (N18, N8, N3, N12);
xor XOR2 (N19, N10, N13);
not NOT1 (N20, N3);
nor NOR2 (N21, N14, N10);
buf BUF1 (N22, N13);
xor XOR2 (N23, N10, N14);
buf BUF1 (N24, N10);
and AND3 (N25, N4, N18, N16);
xor XOR2 (N26, N12, N6);
buf BUF1 (N27, N10);
buf BUF1 (N28, N22);
nor NOR2 (N29, N21, N13);
buf BUF1 (N30, N20);
nor NOR3 (N31, N26, N8, N29);
or OR3 (N32, N3, N16, N15);
xor XOR2 (N33, N26, N17);
buf BUF1 (N34, N25);
and AND3 (N35, N30, N6, N13);
xor XOR2 (N36, N27, N15);
not NOT1 (N37, N28);
xor XOR2 (N38, N34, N20);
not NOT1 (N39, N36);
not NOT1 (N40, N23);
and AND2 (N41, N37, N9);
or OR2 (N42, N24, N2);
not NOT1 (N43, N40);
xor XOR2 (N44, N41, N3);
or OR4 (N45, N32, N6, N10, N15);
nand NAND2 (N46, N44, N27);
xor XOR2 (N47, N19, N33);
nand NAND2 (N48, N27, N27);
nor NOR3 (N49, N39, N25, N22);
and AND2 (N50, N47, N8);
and AND3 (N51, N48, N15, N15);
nor NOR4 (N52, N49, N49, N43, N8);
nor NOR4 (N53, N49, N32, N41, N46);
or OR2 (N54, N28, N35);
not NOT1 (N55, N38);
or OR3 (N56, N8, N28, N53);
or OR4 (N57, N30, N53, N56, N12);
nand NAND3 (N58, N43, N45, N31);
not NOT1 (N59, N7);
nor NOR4 (N60, N39, N13, N53, N42);
nor NOR2 (N61, N30, N19);
xor XOR2 (N62, N59, N8);
buf BUF1 (N63, N50);
or OR3 (N64, N61, N51, N23);
not NOT1 (N65, N46);
nor NOR2 (N66, N65, N26);
xor XOR2 (N67, N64, N5);
not NOT1 (N68, N60);
and AND3 (N69, N52, N65, N40);
xor XOR2 (N70, N55, N13);
or OR4 (N71, N68, N43, N14, N59);
and AND4 (N72, N57, N41, N51, N22);
or OR4 (N73, N67, N4, N58, N8);
not NOT1 (N74, N47);
xor XOR2 (N75, N72, N25);
nand NAND3 (N76, N63, N28, N52);
or OR2 (N77, N62, N43);
or OR4 (N78, N73, N54, N73, N66);
not NOT1 (N79, N36);
buf BUF1 (N80, N21);
xor XOR2 (N81, N79, N30);
or OR3 (N82, N74, N40, N30);
xor XOR2 (N83, N75, N75);
nor NOR3 (N84, N81, N62, N62);
nor NOR2 (N85, N83, N12);
or OR4 (N86, N70, N79, N81, N4);
xor XOR2 (N87, N78, N57);
or OR4 (N88, N84, N62, N50, N13);
xor XOR2 (N89, N86, N68);
xor XOR2 (N90, N82, N64);
xor XOR2 (N91, N88, N80);
buf BUF1 (N92, N29);
or OR3 (N93, N77, N18, N52);
buf BUF1 (N94, N93);
xor XOR2 (N95, N89, N61);
and AND3 (N96, N91, N52, N12);
nor NOR4 (N97, N71, N23, N15, N31);
or OR2 (N98, N96, N83);
not NOT1 (N99, N97);
nor NOR4 (N100, N90, N86, N58, N74);
and AND2 (N101, N76, N54);
and AND3 (N102, N92, N100, N96);
buf BUF1 (N103, N25);
xor XOR2 (N104, N102, N74);
not NOT1 (N105, N95);
xor XOR2 (N106, N69, N2);
xor XOR2 (N107, N98, N11);
or OR4 (N108, N94, N99, N70, N83);
nor NOR3 (N109, N53, N104, N9);
nor NOR3 (N110, N34, N68, N100);
not NOT1 (N111, N87);
xor XOR2 (N112, N108, N63);
not NOT1 (N113, N112);
nand NAND3 (N114, N109, N24, N11);
not NOT1 (N115, N107);
and AND2 (N116, N114, N115);
nor NOR3 (N117, N16, N62, N3);
and AND3 (N118, N113, N104, N86);
buf BUF1 (N119, N103);
not NOT1 (N120, N85);
and AND4 (N121, N110, N54, N42, N109);
buf BUF1 (N122, N106);
or OR2 (N123, N116, N14);
not NOT1 (N124, N118);
nor NOR2 (N125, N123, N54);
or OR4 (N126, N125, N111, N119, N12);
not NOT1 (N127, N19);
xor XOR2 (N128, N121, N65);
nand NAND2 (N129, N24, N79);
buf BUF1 (N130, N129);
buf BUF1 (N131, N130);
nand NAND3 (N132, N117, N97, N25);
buf BUF1 (N133, N105);
nor NOR2 (N134, N127, N53);
nand NAND2 (N135, N120, N8);
not NOT1 (N136, N101);
nor NOR2 (N137, N131, N5);
xor XOR2 (N138, N122, N76);
nor NOR3 (N139, N124, N104, N104);
buf BUF1 (N140, N136);
nor NOR3 (N141, N140, N57, N61);
or OR4 (N142, N139, N47, N113, N137);
or OR2 (N143, N12, N103);
nand NAND3 (N144, N133, N137, N34);
buf BUF1 (N145, N132);
not NOT1 (N146, N142);
nand NAND3 (N147, N138, N6, N59);
not NOT1 (N148, N134);
nor NOR4 (N149, N126, N111, N97, N140);
xor XOR2 (N150, N135, N111);
xor XOR2 (N151, N144, N90);
or OR2 (N152, N151, N87);
nand NAND4 (N153, N146, N87, N128, N61);
or OR4 (N154, N52, N82, N40, N108);
buf BUF1 (N155, N143);
or OR2 (N156, N149, N136);
buf BUF1 (N157, N154);
buf BUF1 (N158, N147);
not NOT1 (N159, N156);
or OR4 (N160, N145, N31, N41, N110);
and AND2 (N161, N153, N142);
buf BUF1 (N162, N159);
not NOT1 (N163, N150);
buf BUF1 (N164, N157);
not NOT1 (N165, N164);
not NOT1 (N166, N152);
and AND2 (N167, N162, N15);
buf BUF1 (N168, N141);
nand NAND3 (N169, N163, N94, N6);
and AND4 (N170, N165, N152, N115, N156);
buf BUF1 (N171, N170);
or OR3 (N172, N148, N11, N116);
not NOT1 (N173, N171);
nor NOR2 (N174, N161, N83);
xor XOR2 (N175, N166, N85);
buf BUF1 (N176, N174);
nand NAND4 (N177, N173, N147, N96, N172);
nand NAND2 (N178, N88, N41);
nand NAND2 (N179, N155, N89);
nor NOR4 (N180, N169, N36, N35, N27);
and AND2 (N181, N180, N81);
not NOT1 (N182, N160);
xor XOR2 (N183, N179, N57);
buf BUF1 (N184, N175);
not NOT1 (N185, N167);
or OR4 (N186, N181, N32, N28, N111);
and AND2 (N187, N182, N42);
or OR2 (N188, N187, N20);
nand NAND3 (N189, N177, N165, N143);
buf BUF1 (N190, N183);
nand NAND4 (N191, N186, N167, N91, N43);
not NOT1 (N192, N185);
not NOT1 (N193, N176);
and AND2 (N194, N189, N61);
nand NAND2 (N195, N168, N96);
not NOT1 (N196, N195);
or OR2 (N197, N192, N139);
or OR2 (N198, N184, N24);
nand NAND4 (N199, N194, N79, N141, N121);
or OR2 (N200, N193, N126);
buf BUF1 (N201, N158);
nand NAND2 (N202, N191, N50);
or OR4 (N203, N178, N101, N144, N64);
or OR2 (N204, N202, N203);
nand NAND2 (N205, N46, N203);
buf BUF1 (N206, N197);
and AND4 (N207, N200, N88, N12, N64);
nand NAND3 (N208, N190, N63, N183);
nand NAND3 (N209, N198, N171, N5);
nor NOR4 (N210, N204, N74, N9, N78);
not NOT1 (N211, N206);
not NOT1 (N212, N199);
xor XOR2 (N213, N205, N31);
buf BUF1 (N214, N196);
not NOT1 (N215, N209);
nand NAND3 (N216, N215, N63, N177);
or OR4 (N217, N207, N169, N215, N91);
nand NAND4 (N218, N208, N75, N36, N99);
nor NOR4 (N219, N212, N153, N81, N93);
nor NOR4 (N220, N219, N162, N101, N26);
or OR4 (N221, N213, N89, N125, N96);
xor XOR2 (N222, N211, N157);
not NOT1 (N223, N217);
buf BUF1 (N224, N216);
or OR4 (N225, N220, N180, N98, N92);
nand NAND2 (N226, N224, N170);
nor NOR2 (N227, N223, N104);
not NOT1 (N228, N210);
nand NAND2 (N229, N225, N25);
nor NOR2 (N230, N188, N82);
buf BUF1 (N231, N228);
xor XOR2 (N232, N214, N58);
nand NAND2 (N233, N221, N202);
not NOT1 (N234, N232);
xor XOR2 (N235, N231, N104);
or OR3 (N236, N234, N65, N67);
xor XOR2 (N237, N222, N183);
nand NAND4 (N238, N229, N208, N228, N88);
buf BUF1 (N239, N238);
not NOT1 (N240, N235);
nor NOR4 (N241, N201, N76, N155, N59);
buf BUF1 (N242, N230);
nand NAND3 (N243, N227, N186, N216);
or OR2 (N244, N236, N120);
nand NAND4 (N245, N241, N57, N42, N116);
nor NOR4 (N246, N242, N176, N90, N13);
buf BUF1 (N247, N240);
and AND2 (N248, N244, N47);
nand NAND2 (N249, N237, N193);
nand NAND3 (N250, N226, N208, N53);
xor XOR2 (N251, N218, N38);
not NOT1 (N252, N239);
not NOT1 (N253, N249);
not NOT1 (N254, N253);
nor NOR2 (N255, N250, N123);
nor NOR2 (N256, N251, N90);
xor XOR2 (N257, N252, N43);
and AND4 (N258, N255, N246, N111, N106);
and AND4 (N259, N230, N13, N99, N193);
buf BUF1 (N260, N233);
nor NOR4 (N261, N247, N224, N78, N216);
nand NAND4 (N262, N260, N27, N58, N52);
or OR4 (N263, N243, N141, N96, N260);
nand NAND2 (N264, N245, N59);
buf BUF1 (N265, N261);
xor XOR2 (N266, N263, N22);
and AND4 (N267, N265, N74, N20, N173);
or OR2 (N268, N259, N82);
nor NOR3 (N269, N268, N11, N208);
buf BUF1 (N270, N257);
or OR2 (N271, N254, N222);
nor NOR2 (N272, N256, N63);
and AND4 (N273, N262, N56, N221, N166);
nand NAND2 (N274, N248, N131);
xor XOR2 (N275, N272, N50);
and AND4 (N276, N258, N230, N152, N83);
nor NOR2 (N277, N276, N275);
and AND2 (N278, N251, N167);
or OR2 (N279, N266, N225);
and AND4 (N280, N270, N108, N81, N162);
not NOT1 (N281, N264);
buf BUF1 (N282, N281);
xor XOR2 (N283, N279, N271);
buf BUF1 (N284, N205);
buf BUF1 (N285, N284);
xor XOR2 (N286, N282, N230);
xor XOR2 (N287, N278, N139);
nand NAND2 (N288, N280, N56);
nand NAND3 (N289, N277, N219, N277);
nand NAND3 (N290, N286, N146, N8);
nand NAND4 (N291, N273, N167, N290, N175);
buf BUF1 (N292, N175);
or OR3 (N293, N292, N44, N180);
not NOT1 (N294, N269);
xor XOR2 (N295, N267, N271);
buf BUF1 (N296, N283);
and AND2 (N297, N289, N68);
nand NAND3 (N298, N297, N254, N56);
nor NOR4 (N299, N291, N268, N293, N33);
nor NOR2 (N300, N199, N110);
or OR2 (N301, N296, N51);
or OR3 (N302, N287, N150, N25);
and AND4 (N303, N299, N125, N225, N145);
not NOT1 (N304, N298);
nor NOR3 (N305, N274, N282, N109);
not NOT1 (N306, N302);
xor XOR2 (N307, N304, N250);
buf BUF1 (N308, N300);
not NOT1 (N309, N308);
xor XOR2 (N310, N295, N297);
nor NOR4 (N311, N305, N290, N233, N38);
nor NOR4 (N312, N294, N18, N195, N113);
and AND4 (N313, N303, N254, N170, N254);
and AND2 (N314, N310, N67);
buf BUF1 (N315, N309);
buf BUF1 (N316, N285);
nor NOR4 (N317, N314, N250, N89, N255);
xor XOR2 (N318, N307, N184);
and AND3 (N319, N312, N9, N48);
or OR2 (N320, N318, N247);
not NOT1 (N321, N301);
and AND3 (N322, N311, N98, N241);
or OR2 (N323, N306, N231);
not NOT1 (N324, N288);
buf BUF1 (N325, N323);
not NOT1 (N326, N319);
buf BUF1 (N327, N320);
and AND3 (N328, N324, N15, N186);
not NOT1 (N329, N321);
xor XOR2 (N330, N322, N122);
buf BUF1 (N331, N315);
not NOT1 (N332, N313);
not NOT1 (N333, N331);
xor XOR2 (N334, N317, N89);
and AND3 (N335, N329, N140, N113);
not NOT1 (N336, N335);
buf BUF1 (N337, N327);
nor NOR3 (N338, N328, N133, N72);
nand NAND2 (N339, N336, N163);
xor XOR2 (N340, N338, N138);
not NOT1 (N341, N334);
and AND2 (N342, N332, N73);
buf BUF1 (N343, N340);
nand NAND4 (N344, N316, N303, N32, N171);
not NOT1 (N345, N341);
and AND3 (N346, N339, N56, N56);
nand NAND3 (N347, N330, N12, N221);
nor NOR3 (N348, N346, N202, N209);
or OR4 (N349, N345, N226, N176, N344);
or OR2 (N350, N247, N278);
nor NOR3 (N351, N348, N303, N219);
nand NAND4 (N352, N342, N335, N42, N231);
nor NOR3 (N353, N333, N21, N188);
xor XOR2 (N354, N349, N167);
and AND2 (N355, N326, N239);
xor XOR2 (N356, N347, N220);
or OR4 (N357, N337, N19, N114, N10);
or OR3 (N358, N350, N81, N249);
buf BUF1 (N359, N356);
nand NAND2 (N360, N354, N2);
not NOT1 (N361, N358);
or OR2 (N362, N359, N150);
or OR4 (N363, N361, N172, N23, N284);
nor NOR3 (N364, N360, N104, N43);
buf BUF1 (N365, N355);
and AND2 (N366, N353, N124);
buf BUF1 (N367, N363);
and AND2 (N368, N325, N335);
nand NAND4 (N369, N362, N353, N5, N129);
not NOT1 (N370, N366);
buf BUF1 (N371, N343);
nand NAND3 (N372, N370, N52, N44);
or OR4 (N373, N367, N44, N370, N65);
not NOT1 (N374, N357);
xor XOR2 (N375, N364, N189);
not NOT1 (N376, N368);
or OR2 (N377, N371, N136);
nand NAND4 (N378, N351, N365, N342, N172);
buf BUF1 (N379, N332);
not NOT1 (N380, N377);
and AND2 (N381, N378, N160);
or OR2 (N382, N375, N234);
nand NAND3 (N383, N380, N209, N239);
not NOT1 (N384, N373);
nor NOR2 (N385, N379, N168);
buf BUF1 (N386, N383);
nand NAND3 (N387, N369, N36, N189);
buf BUF1 (N388, N384);
xor XOR2 (N389, N352, N89);
nor NOR2 (N390, N376, N216);
nor NOR2 (N391, N385, N199);
or OR3 (N392, N389, N14, N16);
and AND4 (N393, N390, N388, N48, N64);
or OR2 (N394, N356, N366);
nor NOR4 (N395, N382, N237, N368, N257);
or OR4 (N396, N391, N322, N298, N167);
not NOT1 (N397, N387);
xor XOR2 (N398, N397, N45);
xor XOR2 (N399, N374, N55);
not NOT1 (N400, N372);
buf BUF1 (N401, N386);
buf BUF1 (N402, N401);
and AND4 (N403, N394, N288, N23, N207);
or OR2 (N404, N403, N300);
or OR4 (N405, N395, N60, N231, N319);
buf BUF1 (N406, N392);
xor XOR2 (N407, N398, N356);
and AND3 (N408, N399, N251, N224);
not NOT1 (N409, N406);
not NOT1 (N410, N396);
buf BUF1 (N411, N407);
buf BUF1 (N412, N408);
nand NAND4 (N413, N400, N277, N389, N261);
buf BUF1 (N414, N393);
or OR2 (N415, N411, N364);
xor XOR2 (N416, N414, N79);
xor XOR2 (N417, N404, N17);
not NOT1 (N418, N409);
nand NAND2 (N419, N410, N284);
xor XOR2 (N420, N413, N374);
not NOT1 (N421, N405);
nand NAND3 (N422, N419, N278, N193);
and AND3 (N423, N402, N122, N401);
buf BUF1 (N424, N421);
buf BUF1 (N425, N412);
not NOT1 (N426, N422);
not NOT1 (N427, N417);
not NOT1 (N428, N416);
or OR4 (N429, N427, N252, N191, N189);
or OR3 (N430, N429, N160, N51);
nor NOR2 (N431, N424, N111);
not NOT1 (N432, N381);
buf BUF1 (N433, N428);
buf BUF1 (N434, N415);
not NOT1 (N435, N423);
xor XOR2 (N436, N418, N70);
and AND2 (N437, N426, N241);
not NOT1 (N438, N431);
nand NAND2 (N439, N435, N308);
not NOT1 (N440, N436);
and AND3 (N441, N425, N177, N28);
not NOT1 (N442, N437);
nand NAND2 (N443, N433, N62);
nor NOR2 (N444, N441, N233);
and AND2 (N445, N420, N22);
buf BUF1 (N446, N434);
buf BUF1 (N447, N445);
buf BUF1 (N448, N439);
or OR4 (N449, N448, N1, N309, N238);
xor XOR2 (N450, N446, N3);
nand NAND3 (N451, N432, N176, N295);
and AND3 (N452, N451, N87, N235);
buf BUF1 (N453, N444);
not NOT1 (N454, N443);
buf BUF1 (N455, N453);
nor NOR2 (N456, N447, N189);
and AND3 (N457, N430, N120, N388);
nor NOR2 (N458, N442, N156);
and AND2 (N459, N457, N237);
nor NOR3 (N460, N454, N1, N90);
buf BUF1 (N461, N450);
xor XOR2 (N462, N456, N229);
buf BUF1 (N463, N460);
xor XOR2 (N464, N438, N88);
nand NAND2 (N465, N461, N357);
xor XOR2 (N466, N464, N33);
buf BUF1 (N467, N459);
not NOT1 (N468, N455);
nand NAND2 (N469, N449, N257);
nand NAND2 (N470, N462, N224);
not NOT1 (N471, N465);
or OR4 (N472, N468, N37, N471, N368);
or OR3 (N473, N257, N418, N291);
not NOT1 (N474, N458);
not NOT1 (N475, N469);
or OR3 (N476, N440, N74, N101);
not NOT1 (N477, N473);
and AND2 (N478, N477, N292);
not NOT1 (N479, N474);
nand NAND4 (N480, N476, N271, N250, N346);
not NOT1 (N481, N480);
buf BUF1 (N482, N475);
or OR2 (N483, N481, N333);
nand NAND4 (N484, N483, N236, N15, N129);
nand NAND4 (N485, N470, N192, N47, N348);
nor NOR3 (N486, N484, N315, N163);
nand NAND2 (N487, N466, N401);
nand NAND2 (N488, N487, N247);
buf BUF1 (N489, N467);
xor XOR2 (N490, N488, N381);
nand NAND3 (N491, N485, N327, N119);
and AND2 (N492, N479, N75);
xor XOR2 (N493, N491, N2);
xor XOR2 (N494, N486, N439);
and AND2 (N495, N489, N470);
xor XOR2 (N496, N492, N434);
not NOT1 (N497, N490);
buf BUF1 (N498, N472);
and AND4 (N499, N498, N218, N373, N40);
nand NAND3 (N500, N452, N164, N198);
and AND2 (N501, N493, N150);
nand NAND4 (N502, N478, N162, N255, N212);
xor XOR2 (N503, N497, N295);
xor XOR2 (N504, N499, N253);
and AND3 (N505, N482, N219, N384);
nand NAND3 (N506, N496, N472, N395);
xor XOR2 (N507, N495, N255);
and AND3 (N508, N494, N187, N58);
buf BUF1 (N509, N508);
not NOT1 (N510, N463);
nand NAND4 (N511, N506, N276, N310, N16);
nand NAND2 (N512, N505, N89);
nor NOR3 (N513, N500, N54, N282);
xor XOR2 (N514, N507, N376);
not NOT1 (N515, N514);
nand NAND2 (N516, N503, N340);
nor NOR4 (N517, N509, N162, N139, N246);
nand NAND4 (N518, N515, N272, N363, N339);
nor NOR2 (N519, N517, N456);
nor NOR3 (N520, N504, N323, N325);
and AND4 (N521, N510, N477, N167, N43);
buf BUF1 (N522, N516);
and AND4 (N523, N520, N458, N146, N237);
nand NAND3 (N524, N523, N189, N71);
and AND2 (N525, N511, N109);
or OR2 (N526, N525, N297);
and AND4 (N527, N521, N72, N199, N462);
and AND4 (N528, N513, N314, N49, N196);
nor NOR3 (N529, N518, N234, N82);
not NOT1 (N530, N519);
nand NAND3 (N531, N522, N306, N259);
nor NOR2 (N532, N529, N215);
nor NOR4 (N533, N526, N331, N359, N354);
not NOT1 (N534, N524);
xor XOR2 (N535, N501, N321);
buf BUF1 (N536, N512);
nand NAND2 (N537, N530, N254);
not NOT1 (N538, N527);
and AND4 (N539, N535, N259, N279, N195);
not NOT1 (N540, N531);
nand NAND2 (N541, N539, N423);
and AND2 (N542, N502, N506);
xor XOR2 (N543, N533, N332);
and AND4 (N544, N538, N486, N33, N307);
nor NOR2 (N545, N541, N136);
and AND2 (N546, N540, N308);
nand NAND3 (N547, N532, N192, N237);
buf BUF1 (N548, N528);
nor NOR3 (N549, N548, N322, N11);
buf BUF1 (N550, N545);
xor XOR2 (N551, N549, N431);
or OR3 (N552, N547, N173, N380);
not NOT1 (N553, N544);
and AND2 (N554, N542, N418);
nor NOR2 (N555, N536, N535);
nand NAND3 (N556, N553, N99, N271);
and AND4 (N557, N550, N147, N130, N442);
or OR3 (N558, N551, N85, N159);
nand NAND2 (N559, N537, N481);
or OR2 (N560, N557, N503);
nand NAND4 (N561, N543, N435, N150, N354);
or OR2 (N562, N534, N407);
and AND3 (N563, N555, N204, N484);
nor NOR4 (N564, N561, N382, N317, N113);
xor XOR2 (N565, N560, N324);
nor NOR2 (N566, N558, N29);
and AND3 (N567, N562, N42, N479);
buf BUF1 (N568, N546);
xor XOR2 (N569, N566, N532);
nor NOR2 (N570, N563, N156);
nand NAND2 (N571, N569, N403);
and AND4 (N572, N568, N565, N83, N302);
or OR3 (N573, N157, N307, N446);
buf BUF1 (N574, N559);
xor XOR2 (N575, N567, N222);
nor NOR4 (N576, N573, N72, N337, N499);
and AND2 (N577, N564, N34);
buf BUF1 (N578, N576);
nor NOR2 (N579, N571, N60);
buf BUF1 (N580, N578);
not NOT1 (N581, N572);
and AND3 (N582, N579, N244, N379);
nand NAND3 (N583, N582, N305, N485);
buf BUF1 (N584, N570);
xor XOR2 (N585, N552, N408);
or OR2 (N586, N556, N9);
and AND3 (N587, N586, N480, N154);
or OR4 (N588, N575, N550, N245, N37);
nor NOR2 (N589, N581, N21);
nand NAND4 (N590, N587, N471, N74, N355);
not NOT1 (N591, N589);
or OR4 (N592, N580, N69, N381, N376);
and AND4 (N593, N592, N579, N235, N166);
or OR2 (N594, N577, N435);
xor XOR2 (N595, N554, N18);
buf BUF1 (N596, N594);
nand NAND3 (N597, N584, N350, N594);
or OR4 (N598, N596, N546, N339, N75);
buf BUF1 (N599, N583);
xor XOR2 (N600, N595, N116);
nand NAND2 (N601, N599, N209);
buf BUF1 (N602, N600);
and AND2 (N603, N601, N460);
xor XOR2 (N604, N597, N532);
or OR2 (N605, N602, N143);
not NOT1 (N606, N598);
or OR2 (N607, N591, N235);
buf BUF1 (N608, N585);
not NOT1 (N609, N593);
nand NAND3 (N610, N588, N31, N258);
and AND3 (N611, N603, N544, N262);
nand NAND3 (N612, N607, N415, N512);
nand NAND3 (N613, N574, N35, N172);
nor NOR2 (N614, N590, N102);
and AND2 (N615, N614, N397);
not NOT1 (N616, N611);
or OR4 (N617, N616, N64, N211, N514);
nor NOR2 (N618, N605, N29);
not NOT1 (N619, N612);
not NOT1 (N620, N613);
not NOT1 (N621, N610);
buf BUF1 (N622, N617);
not NOT1 (N623, N618);
buf BUF1 (N624, N609);
not NOT1 (N625, N620);
nor NOR4 (N626, N623, N559, N65, N14);
not NOT1 (N627, N621);
nor NOR4 (N628, N626, N471, N430, N449);
nor NOR4 (N629, N624, N58, N26, N368);
and AND2 (N630, N629, N287);
or OR3 (N631, N628, N544, N377);
and AND3 (N632, N608, N609, N478);
nand NAND4 (N633, N630, N123, N579, N463);
not NOT1 (N634, N627);
buf BUF1 (N635, N606);
buf BUF1 (N636, N635);
nand NAND4 (N637, N604, N227, N312, N62);
and AND2 (N638, N632, N135);
nand NAND3 (N639, N631, N273, N602);
not NOT1 (N640, N625);
or OR3 (N641, N634, N620, N406);
and AND4 (N642, N619, N558, N600, N104);
xor XOR2 (N643, N615, N544);
buf BUF1 (N644, N640);
xor XOR2 (N645, N644, N60);
or OR3 (N646, N636, N550, N150);
or OR4 (N647, N633, N247, N560, N464);
nor NOR2 (N648, N646, N342);
not NOT1 (N649, N637);
not NOT1 (N650, N643);
nor NOR3 (N651, N639, N109, N482);
and AND3 (N652, N641, N152, N226);
nand NAND4 (N653, N642, N243, N514, N49);
xor XOR2 (N654, N645, N601);
xor XOR2 (N655, N649, N372);
nand NAND4 (N656, N638, N651, N407, N445);
nor NOR4 (N657, N33, N11, N542, N625);
nor NOR2 (N658, N622, N255);
or OR3 (N659, N656, N137, N115);
nand NAND4 (N660, N648, N413, N31, N227);
and AND2 (N661, N655, N430);
and AND2 (N662, N659, N55);
nand NAND4 (N663, N658, N158, N556, N8);
nand NAND2 (N664, N652, N152);
or OR2 (N665, N660, N185);
buf BUF1 (N666, N661);
and AND4 (N667, N663, N194, N627, N454);
nand NAND3 (N668, N667, N501, N347);
or OR4 (N669, N665, N117, N341, N161);
nor NOR2 (N670, N647, N270);
and AND2 (N671, N670, N368);
nor NOR2 (N672, N669, N615);
nand NAND3 (N673, N671, N295, N272);
nand NAND2 (N674, N664, N659);
nor NOR2 (N675, N674, N460);
not NOT1 (N676, N657);
and AND3 (N677, N650, N67, N157);
buf BUF1 (N678, N668);
nand NAND3 (N679, N673, N541, N141);
or OR3 (N680, N654, N484, N255);
not NOT1 (N681, N662);
nand NAND3 (N682, N676, N297, N40);
buf BUF1 (N683, N672);
or OR2 (N684, N682, N1);
or OR2 (N685, N679, N423);
not NOT1 (N686, N680);
and AND4 (N687, N683, N123, N52, N133);
xor XOR2 (N688, N681, N603);
nand NAND4 (N689, N678, N289, N267, N479);
nand NAND3 (N690, N686, N194, N84);
and AND3 (N691, N689, N212, N460);
not NOT1 (N692, N653);
not NOT1 (N693, N685);
or OR2 (N694, N691, N53);
xor XOR2 (N695, N677, N130);
xor XOR2 (N696, N695, N17);
xor XOR2 (N697, N692, N285);
and AND4 (N698, N687, N44, N382, N552);
nor NOR3 (N699, N698, N352, N494);
nor NOR4 (N700, N688, N616, N78, N664);
xor XOR2 (N701, N699, N579);
nand NAND3 (N702, N700, N218, N156);
xor XOR2 (N703, N693, N395);
buf BUF1 (N704, N703);
xor XOR2 (N705, N704, N359);
buf BUF1 (N706, N697);
buf BUF1 (N707, N706);
or OR2 (N708, N666, N440);
and AND3 (N709, N684, N694, N221);
and AND4 (N710, N546, N266, N58, N72);
or OR3 (N711, N701, N242, N485);
nor NOR4 (N712, N710, N19, N458, N632);
xor XOR2 (N713, N708, N578);
or OR4 (N714, N675, N12, N357, N697);
nand NAND4 (N715, N712, N521, N110, N2);
and AND3 (N716, N705, N496, N64);
nand NAND2 (N717, N711, N697);
nor NOR2 (N718, N696, N251);
nor NOR4 (N719, N717, N35, N545, N39);
and AND2 (N720, N690, N453);
nand NAND2 (N721, N715, N91);
xor XOR2 (N722, N718, N143);
buf BUF1 (N723, N716);
nor NOR3 (N724, N709, N126, N607);
and AND4 (N725, N722, N605, N403, N245);
xor XOR2 (N726, N723, N591);
and AND3 (N727, N725, N351, N259);
and AND2 (N728, N727, N522);
not NOT1 (N729, N714);
buf BUF1 (N730, N729);
and AND4 (N731, N726, N175, N74, N370);
xor XOR2 (N732, N713, N170);
xor XOR2 (N733, N728, N239);
buf BUF1 (N734, N732);
and AND4 (N735, N733, N63, N215, N235);
buf BUF1 (N736, N720);
buf BUF1 (N737, N734);
buf BUF1 (N738, N735);
nor NOR4 (N739, N702, N310, N312, N5);
or OR3 (N740, N739, N375, N433);
not NOT1 (N741, N707);
and AND4 (N742, N740, N332, N39, N130);
and AND4 (N743, N721, N153, N319, N136);
and AND3 (N744, N724, N281, N58);
nand NAND3 (N745, N731, N17, N128);
nand NAND2 (N746, N745, N724);
not NOT1 (N747, N736);
nand NAND2 (N748, N743, N657);
not NOT1 (N749, N748);
xor XOR2 (N750, N749, N272);
nor NOR2 (N751, N730, N590);
not NOT1 (N752, N738);
nor NOR2 (N753, N750, N561);
nand NAND3 (N754, N747, N611, N8);
xor XOR2 (N755, N754, N726);
nand NAND4 (N756, N751, N84, N542, N77);
and AND2 (N757, N737, N552);
buf BUF1 (N758, N755);
buf BUF1 (N759, N753);
nand NAND2 (N760, N741, N44);
not NOT1 (N761, N719);
buf BUF1 (N762, N757);
nand NAND2 (N763, N744, N719);
or OR4 (N764, N763, N26, N397, N558);
and AND2 (N765, N742, N258);
nor NOR4 (N766, N752, N479, N643, N470);
and AND3 (N767, N766, N458, N631);
nor NOR3 (N768, N756, N501, N750);
nand NAND4 (N769, N764, N138, N391, N343);
and AND4 (N770, N759, N11, N419, N282);
xor XOR2 (N771, N761, N1);
xor XOR2 (N772, N770, N587);
nand NAND4 (N773, N771, N263, N495, N613);
not NOT1 (N774, N760);
buf BUF1 (N775, N768);
not NOT1 (N776, N762);
not NOT1 (N777, N765);
or OR3 (N778, N769, N303, N499);
not NOT1 (N779, N776);
nand NAND3 (N780, N779, N321, N633);
not NOT1 (N781, N772);
buf BUF1 (N782, N774);
not NOT1 (N783, N758);
nor NOR4 (N784, N775, N356, N62, N586);
xor XOR2 (N785, N782, N707);
xor XOR2 (N786, N773, N638);
nand NAND3 (N787, N777, N519, N12);
nand NAND2 (N788, N778, N547);
xor XOR2 (N789, N784, N644);
and AND3 (N790, N783, N556, N629);
or OR2 (N791, N780, N515);
xor XOR2 (N792, N785, N329);
and AND3 (N793, N791, N163, N112);
xor XOR2 (N794, N767, N375);
nand NAND2 (N795, N789, N201);
buf BUF1 (N796, N792);
xor XOR2 (N797, N796, N151);
xor XOR2 (N798, N790, N636);
xor XOR2 (N799, N787, N330);
or OR2 (N800, N797, N647);
xor XOR2 (N801, N799, N211);
not NOT1 (N802, N794);
nor NOR3 (N803, N802, N616, N155);
or OR4 (N804, N793, N80, N193, N696);
and AND3 (N805, N798, N675, N51);
and AND3 (N806, N746, N524, N779);
and AND3 (N807, N781, N45, N290);
nand NAND2 (N808, N795, N412);
not NOT1 (N809, N805);
nor NOR2 (N810, N804, N727);
xor XOR2 (N811, N806, N449);
buf BUF1 (N812, N807);
nor NOR4 (N813, N800, N487, N314, N474);
and AND3 (N814, N813, N172, N123);
and AND4 (N815, N786, N737, N276, N85);
or OR2 (N816, N812, N20);
or OR4 (N817, N811, N816, N26, N699);
buf BUF1 (N818, N488);
nand NAND4 (N819, N815, N200, N585, N141);
nor NOR2 (N820, N818, N20);
nand NAND2 (N821, N817, N66);
nand NAND3 (N822, N814, N622, N186);
xor XOR2 (N823, N820, N725);
not NOT1 (N824, N823);
xor XOR2 (N825, N810, N375);
and AND4 (N826, N821, N309, N428, N108);
not NOT1 (N827, N803);
and AND2 (N828, N819, N225);
or OR2 (N829, N788, N62);
buf BUF1 (N830, N827);
and AND4 (N831, N825, N419, N583, N582);
nor NOR4 (N832, N801, N306, N758, N761);
xor XOR2 (N833, N826, N789);
xor XOR2 (N834, N828, N112);
or OR4 (N835, N834, N804, N251, N106);
buf BUF1 (N836, N808);
and AND2 (N837, N829, N342);
not NOT1 (N838, N809);
buf BUF1 (N839, N835);
not NOT1 (N840, N824);
or OR4 (N841, N832, N245, N122, N501);
nor NOR3 (N842, N822, N551, N313);
not NOT1 (N843, N838);
not NOT1 (N844, N841);
or OR4 (N845, N830, N617, N122, N631);
not NOT1 (N846, N844);
nand NAND4 (N847, N843, N693, N590, N347);
nand NAND2 (N848, N845, N303);
buf BUF1 (N849, N833);
or OR4 (N850, N839, N510, N384, N406);
buf BUF1 (N851, N840);
and AND3 (N852, N847, N680, N55);
nor NOR4 (N853, N846, N564, N200, N388);
and AND2 (N854, N848, N684);
not NOT1 (N855, N849);
not NOT1 (N856, N852);
nor NOR4 (N857, N836, N254, N501, N825);
nand NAND4 (N858, N850, N206, N785, N262);
nor NOR3 (N859, N853, N522, N346);
xor XOR2 (N860, N858, N195);
nor NOR3 (N861, N831, N859, N115);
nand NAND2 (N862, N568, N344);
buf BUF1 (N863, N855);
buf BUF1 (N864, N862);
or OR2 (N865, N863, N547);
nor NOR2 (N866, N837, N159);
and AND2 (N867, N857, N46);
nor NOR3 (N868, N865, N324, N284);
xor XOR2 (N869, N842, N288);
buf BUF1 (N870, N866);
buf BUF1 (N871, N867);
or OR3 (N872, N870, N574, N746);
or OR2 (N873, N869, N853);
xor XOR2 (N874, N864, N557);
xor XOR2 (N875, N868, N822);
xor XOR2 (N876, N856, N814);
nor NOR4 (N877, N875, N663, N113, N141);
not NOT1 (N878, N876);
not NOT1 (N879, N854);
or OR2 (N880, N874, N146);
xor XOR2 (N881, N860, N68);
nand NAND2 (N882, N861, N20);
nor NOR4 (N883, N878, N27, N615, N336);
buf BUF1 (N884, N877);
not NOT1 (N885, N873);
xor XOR2 (N886, N851, N444);
or OR2 (N887, N881, N734);
or OR4 (N888, N885, N599, N493, N324);
nand NAND2 (N889, N882, N653);
or OR3 (N890, N889, N873, N548);
or OR4 (N891, N872, N244, N842, N295);
or OR3 (N892, N884, N609, N380);
xor XOR2 (N893, N879, N833);
not NOT1 (N894, N890);
xor XOR2 (N895, N892, N759);
not NOT1 (N896, N893);
not NOT1 (N897, N887);
nor NOR4 (N898, N896, N21, N224, N165);
nand NAND4 (N899, N886, N37, N797, N593);
or OR3 (N900, N899, N258, N351);
and AND2 (N901, N883, N307);
or OR3 (N902, N895, N829, N427);
and AND2 (N903, N894, N117);
and AND4 (N904, N880, N371, N403, N256);
buf BUF1 (N905, N891);
or OR4 (N906, N898, N729, N411, N66);
xor XOR2 (N907, N904, N236);
nor NOR4 (N908, N871, N175, N267, N455);
not NOT1 (N909, N905);
xor XOR2 (N910, N909, N242);
not NOT1 (N911, N906);
buf BUF1 (N912, N908);
buf BUF1 (N913, N912);
or OR3 (N914, N911, N235, N572);
nor NOR3 (N915, N907, N59, N433);
xor XOR2 (N916, N901, N886);
buf BUF1 (N917, N902);
endmodule