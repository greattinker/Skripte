// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13;

output N2481,N2503,N2478,N2508,N2496,N2499,N2512,N2510,N2500,N2513;

buf BUF1 (N14, N2);
nand NAND3 (N15, N11, N5, N12);
xor XOR2 (N16, N10, N5);
nand NAND4 (N17, N5, N14, N3, N11);
or OR2 (N18, N12, N4);
buf BUF1 (N19, N3);
nor NOR3 (N20, N9, N13, N2);
xor XOR2 (N21, N9, N5);
nor NOR2 (N22, N15, N15);
nor NOR2 (N23, N6, N6);
or OR2 (N24, N16, N14);
nor NOR4 (N25, N22, N8, N17, N19);
and AND4 (N26, N6, N10, N18, N19);
nor NOR3 (N27, N13, N14, N26);
nor NOR3 (N28, N5, N14, N7);
not NOT1 (N29, N20);
not NOT1 (N30, N12);
and AND4 (N31, N18, N14, N6, N13);
buf BUF1 (N32, N14);
and AND4 (N33, N27, N8, N32, N12);
xor XOR2 (N34, N29, N17);
nor NOR4 (N35, N14, N13, N31, N19);
not NOT1 (N36, N9);
and AND4 (N37, N28, N4, N33, N5);
buf BUF1 (N38, N33);
buf BUF1 (N39, N34);
or OR3 (N40, N37, N15, N29);
nand NAND4 (N41, N35, N2, N40, N39);
xor XOR2 (N42, N37, N22);
nand NAND2 (N43, N39, N14);
not NOT1 (N44, N30);
nor NOR3 (N45, N21, N20, N34);
or OR2 (N46, N44, N30);
buf BUF1 (N47, N36);
or OR2 (N48, N42, N22);
or OR4 (N49, N43, N5, N29, N14);
or OR2 (N50, N25, N39);
buf BUF1 (N51, N47);
not NOT1 (N52, N48);
xor XOR2 (N53, N23, N17);
and AND2 (N54, N52, N18);
xor XOR2 (N55, N45, N47);
buf BUF1 (N56, N24);
or OR2 (N57, N46, N7);
or OR4 (N58, N49, N37, N26, N46);
nand NAND3 (N59, N56, N48, N51);
not NOT1 (N60, N59);
nor NOR4 (N61, N53, N49, N46, N20);
not NOT1 (N62, N30);
not NOT1 (N63, N62);
not NOT1 (N64, N55);
nand NAND3 (N65, N63, N27, N31);
nor NOR4 (N66, N38, N29, N19, N27);
not NOT1 (N67, N66);
not NOT1 (N68, N58);
nor NOR3 (N69, N54, N35, N29);
or OR4 (N70, N67, N28, N26, N36);
nand NAND2 (N71, N61, N69);
nor NOR4 (N72, N63, N15, N49, N41);
nor NOR4 (N73, N11, N14, N46, N44);
xor XOR2 (N74, N71, N21);
and AND2 (N75, N73, N24);
nand NAND3 (N76, N70, N17, N42);
nor NOR2 (N77, N65, N44);
and AND2 (N78, N76, N32);
nor NOR4 (N79, N60, N1, N43, N52);
buf BUF1 (N80, N74);
and AND3 (N81, N57, N59, N70);
not NOT1 (N82, N75);
nand NAND3 (N83, N50, N49, N69);
xor XOR2 (N84, N78, N76);
or OR2 (N85, N81, N15);
not NOT1 (N86, N79);
xor XOR2 (N87, N68, N39);
and AND3 (N88, N85, N57, N48);
xor XOR2 (N89, N87, N62);
not NOT1 (N90, N89);
buf BUF1 (N91, N83);
or OR4 (N92, N82, N53, N71, N77);
nor NOR2 (N93, N33, N54);
buf BUF1 (N94, N86);
and AND4 (N95, N80, N90, N33, N61);
nor NOR3 (N96, N40, N18, N64);
buf BUF1 (N97, N24);
or OR2 (N98, N91, N24);
nor NOR4 (N99, N95, N68, N32, N64);
xor XOR2 (N100, N72, N24);
nand NAND4 (N101, N92, N47, N78, N62);
buf BUF1 (N102, N94);
and AND2 (N103, N93, N8);
not NOT1 (N104, N96);
nor NOR4 (N105, N101, N26, N19, N24);
or OR3 (N106, N102, N51, N97);
and AND2 (N107, N103, N82);
buf BUF1 (N108, N67);
buf BUF1 (N109, N88);
buf BUF1 (N110, N106);
not NOT1 (N111, N105);
buf BUF1 (N112, N111);
and AND2 (N113, N110, N35);
nor NOR3 (N114, N113, N31, N43);
nand NAND2 (N115, N112, N24);
nor NOR3 (N116, N84, N75, N75);
buf BUF1 (N117, N104);
not NOT1 (N118, N107);
nand NAND3 (N119, N99, N5, N31);
xor XOR2 (N120, N109, N25);
not NOT1 (N121, N108);
and AND4 (N122, N98, N70, N103, N57);
nand NAND2 (N123, N119, N109);
nand NAND4 (N124, N114, N3, N82, N2);
and AND2 (N125, N117, N27);
not NOT1 (N126, N121);
and AND2 (N127, N122, N125);
not NOT1 (N128, N33);
and AND2 (N129, N124, N100);
and AND3 (N130, N91, N4, N128);
and AND4 (N131, N73, N104, N31, N97);
buf BUF1 (N132, N127);
or OR4 (N133, N132, N18, N1, N99);
and AND2 (N134, N133, N76);
not NOT1 (N135, N126);
and AND2 (N136, N134, N7);
buf BUF1 (N137, N130);
or OR3 (N138, N115, N63, N17);
nor NOR4 (N139, N129, N93, N127, N38);
xor XOR2 (N140, N123, N36);
and AND4 (N141, N136, N62, N93, N92);
buf BUF1 (N142, N140);
xor XOR2 (N143, N142, N49);
and AND2 (N144, N137, N124);
or OR3 (N145, N120, N49, N42);
not NOT1 (N146, N116);
xor XOR2 (N147, N139, N71);
or OR4 (N148, N118, N138, N2, N48);
and AND3 (N149, N100, N21, N139);
xor XOR2 (N150, N131, N81);
nand NAND4 (N151, N147, N86, N1, N109);
or OR2 (N152, N148, N127);
xor XOR2 (N153, N150, N23);
not NOT1 (N154, N141);
nor NOR4 (N155, N154, N10, N26, N141);
buf BUF1 (N156, N155);
and AND3 (N157, N151, N71, N151);
or OR4 (N158, N156, N136, N82, N21);
not NOT1 (N159, N157);
and AND2 (N160, N135, N109);
nor NOR4 (N161, N143, N10, N21, N38);
xor XOR2 (N162, N159, N117);
xor XOR2 (N163, N158, N100);
not NOT1 (N164, N146);
and AND4 (N165, N153, N87, N145, N9);
or OR2 (N166, N161, N54);
nor NOR2 (N167, N98, N42);
xor XOR2 (N168, N164, N102);
or OR3 (N169, N165, N130, N15);
buf BUF1 (N170, N160);
and AND4 (N171, N162, N35, N73, N96);
nand NAND3 (N172, N152, N139, N139);
and AND3 (N173, N167, N72, N148);
not NOT1 (N174, N149);
nand NAND4 (N175, N166, N72, N137, N23);
xor XOR2 (N176, N173, N102);
nor NOR4 (N177, N172, N139, N70, N112);
and AND4 (N178, N174, N138, N85, N9);
buf BUF1 (N179, N175);
xor XOR2 (N180, N179, N51);
and AND2 (N181, N170, N121);
nor NOR2 (N182, N176, N167);
nand NAND3 (N183, N177, N59, N100);
and AND4 (N184, N169, N182, N10, N57);
buf BUF1 (N185, N19);
nor NOR3 (N186, N178, N34, N179);
nand NAND3 (N187, N183, N57, N80);
xor XOR2 (N188, N163, N140);
or OR3 (N189, N185, N157, N114);
not NOT1 (N190, N186);
nand NAND4 (N191, N168, N67, N182, N83);
buf BUF1 (N192, N181);
nor NOR3 (N193, N180, N24, N123);
not NOT1 (N194, N192);
buf BUF1 (N195, N191);
xor XOR2 (N196, N188, N146);
not NOT1 (N197, N194);
buf BUF1 (N198, N196);
nor NOR2 (N199, N193, N106);
not NOT1 (N200, N190);
not NOT1 (N201, N199);
not NOT1 (N202, N197);
and AND2 (N203, N201, N181);
not NOT1 (N204, N144);
or OR2 (N205, N204, N160);
not NOT1 (N206, N205);
and AND2 (N207, N202, N204);
nor NOR4 (N208, N187, N206, N30, N138);
nor NOR3 (N209, N75, N80, N79);
or OR2 (N210, N195, N132);
or OR2 (N211, N198, N175);
or OR2 (N212, N189, N43);
or OR2 (N213, N212, N4);
xor XOR2 (N214, N208, N81);
buf BUF1 (N215, N200);
and AND2 (N216, N209, N176);
not NOT1 (N217, N216);
buf BUF1 (N218, N213);
nand NAND2 (N219, N211, N195);
xor XOR2 (N220, N219, N147);
and AND2 (N221, N217, N94);
nand NAND3 (N222, N221, N197, N71);
or OR4 (N223, N171, N74, N202, N27);
nor NOR3 (N224, N215, N212, N66);
xor XOR2 (N225, N214, N56);
buf BUF1 (N226, N222);
xor XOR2 (N227, N210, N171);
or OR3 (N228, N226, N141, N120);
nor NOR4 (N229, N224, N103, N191, N34);
nor NOR4 (N230, N225, N47, N115, N182);
buf BUF1 (N231, N228);
nand NAND3 (N232, N184, N107, N158);
and AND2 (N233, N203, N60);
nor NOR4 (N234, N233, N125, N48, N139);
and AND4 (N235, N230, N99, N63, N31);
nor NOR3 (N236, N234, N145, N91);
nand NAND4 (N237, N229, N125, N195, N2);
nor NOR2 (N238, N223, N173);
nor NOR4 (N239, N207, N209, N160, N37);
buf BUF1 (N240, N231);
not NOT1 (N241, N235);
nor NOR4 (N242, N232, N201, N116, N39);
or OR4 (N243, N241, N4, N220, N177);
nand NAND4 (N244, N84, N230, N232, N99);
nand NAND4 (N245, N238, N42, N163, N132);
and AND2 (N246, N242, N122);
nand NAND4 (N247, N236, N199, N132, N57);
xor XOR2 (N248, N245, N244);
or OR2 (N249, N118, N167);
not NOT1 (N250, N239);
or OR4 (N251, N250, N73, N62, N136);
nand NAND3 (N252, N248, N13, N213);
and AND3 (N253, N252, N167, N177);
nand NAND4 (N254, N246, N242, N248, N35);
not NOT1 (N255, N243);
or OR4 (N256, N237, N39, N62, N47);
nor NOR4 (N257, N255, N132, N22, N252);
not NOT1 (N258, N254);
not NOT1 (N259, N240);
xor XOR2 (N260, N227, N19);
xor XOR2 (N261, N218, N120);
or OR4 (N262, N256, N70, N83, N112);
nor NOR4 (N263, N262, N168, N217, N21);
xor XOR2 (N264, N247, N88);
nand NAND4 (N265, N253, N236, N133, N133);
nand NAND3 (N266, N261, N129, N2);
not NOT1 (N267, N265);
buf BUF1 (N268, N249);
buf BUF1 (N269, N258);
and AND3 (N270, N257, N136, N165);
xor XOR2 (N271, N264, N130);
buf BUF1 (N272, N260);
not NOT1 (N273, N266);
nand NAND2 (N274, N267, N260);
xor XOR2 (N275, N263, N269);
nand NAND2 (N276, N70, N144);
xor XOR2 (N277, N259, N93);
xor XOR2 (N278, N270, N160);
buf BUF1 (N279, N271);
buf BUF1 (N280, N268);
xor XOR2 (N281, N273, N236);
and AND4 (N282, N277, N186, N121, N176);
or OR4 (N283, N281, N93, N98, N90);
xor XOR2 (N284, N280, N187);
not NOT1 (N285, N275);
xor XOR2 (N286, N274, N180);
nor NOR4 (N287, N276, N242, N249, N93);
not NOT1 (N288, N272);
xor XOR2 (N289, N286, N182);
and AND3 (N290, N282, N156, N120);
or OR2 (N291, N278, N215);
nand NAND2 (N292, N288, N121);
xor XOR2 (N293, N279, N283);
or OR4 (N294, N194, N7, N151, N240);
not NOT1 (N295, N284);
nand NAND4 (N296, N290, N52, N255, N197);
or OR2 (N297, N289, N95);
and AND4 (N298, N294, N255, N147, N284);
nor NOR4 (N299, N295, N81, N223, N116);
xor XOR2 (N300, N285, N65);
nor NOR2 (N301, N296, N58);
and AND4 (N302, N251, N39, N59, N172);
nand NAND2 (N303, N300, N278);
xor XOR2 (N304, N297, N248);
or OR2 (N305, N291, N84);
not NOT1 (N306, N303);
or OR3 (N307, N305, N229, N38);
nand NAND4 (N308, N299, N26, N219, N232);
buf BUF1 (N309, N304);
buf BUF1 (N310, N307);
and AND2 (N311, N310, N134);
nand NAND2 (N312, N298, N183);
and AND4 (N313, N311, N239, N281, N119);
not NOT1 (N314, N292);
xor XOR2 (N315, N314, N77);
or OR3 (N316, N293, N34, N297);
not NOT1 (N317, N312);
and AND4 (N318, N301, N112, N20, N11);
nor NOR3 (N319, N315, N299, N7);
not NOT1 (N320, N308);
nand NAND4 (N321, N309, N88, N24, N60);
and AND4 (N322, N318, N77, N170, N113);
nand NAND2 (N323, N317, N155);
nand NAND4 (N324, N319, N166, N122, N30);
nand NAND3 (N325, N287, N119, N4);
or OR3 (N326, N320, N193, N315);
not NOT1 (N327, N302);
nor NOR3 (N328, N313, N187, N136);
nand NAND4 (N329, N325, N142, N75, N38);
buf BUF1 (N330, N327);
not NOT1 (N331, N323);
buf BUF1 (N332, N328);
not NOT1 (N333, N306);
nor NOR4 (N334, N329, N173, N15, N182);
not NOT1 (N335, N326);
xor XOR2 (N336, N322, N132);
xor XOR2 (N337, N330, N72);
or OR2 (N338, N337, N146);
and AND2 (N339, N338, N62);
xor XOR2 (N340, N339, N20);
not NOT1 (N341, N331);
and AND2 (N342, N321, N103);
and AND3 (N343, N324, N118, N148);
nand NAND2 (N344, N332, N296);
nand NAND3 (N345, N344, N35, N273);
nand NAND2 (N346, N340, N61);
nand NAND4 (N347, N341, N194, N186, N299);
nor NOR2 (N348, N334, N20);
nand NAND4 (N349, N345, N237, N94, N196);
nor NOR3 (N350, N336, N325, N321);
or OR4 (N351, N349, N39, N282, N265);
and AND3 (N352, N351, N51, N341);
buf BUF1 (N353, N333);
nand NAND4 (N354, N343, N70, N351, N157);
or OR3 (N355, N316, N271, N60);
xor XOR2 (N356, N352, N176);
not NOT1 (N357, N346);
nor NOR4 (N358, N335, N215, N262, N19);
or OR4 (N359, N357, N299, N194, N235);
and AND2 (N360, N350, N207);
nor NOR4 (N361, N348, N83, N225, N235);
or OR4 (N362, N356, N218, N162, N224);
and AND3 (N363, N361, N84, N80);
and AND4 (N364, N359, N129, N33, N363);
nor NOR4 (N365, N315, N167, N265, N214);
not NOT1 (N366, N342);
or OR4 (N367, N358, N224, N253, N87);
nor NOR4 (N368, N362, N31, N104, N298);
buf BUF1 (N369, N353);
nor NOR2 (N370, N364, N202);
nor NOR4 (N371, N367, N222, N21, N194);
and AND3 (N372, N371, N266, N160);
nor NOR4 (N373, N372, N66, N147, N145);
nand NAND3 (N374, N355, N162, N216);
and AND2 (N375, N365, N359);
xor XOR2 (N376, N369, N222);
and AND4 (N377, N373, N50, N158, N346);
or OR3 (N378, N370, N241, N246);
or OR4 (N379, N368, N28, N156, N260);
or OR3 (N380, N378, N108, N14);
nand NAND2 (N381, N366, N190);
xor XOR2 (N382, N379, N143);
and AND4 (N383, N376, N261, N237, N364);
nand NAND2 (N384, N354, N41);
and AND3 (N385, N374, N170, N44);
nor NOR2 (N386, N377, N362);
not NOT1 (N387, N380);
buf BUF1 (N388, N382);
buf BUF1 (N389, N360);
and AND3 (N390, N383, N260, N11);
xor XOR2 (N391, N387, N387);
or OR4 (N392, N384, N349, N390, N3);
nand NAND3 (N393, N309, N72, N60);
buf BUF1 (N394, N381);
nor NOR2 (N395, N391, N155);
or OR2 (N396, N388, N369);
or OR3 (N397, N386, N151, N251);
xor XOR2 (N398, N347, N246);
nand NAND3 (N399, N375, N13, N162);
and AND3 (N400, N398, N112, N5);
and AND3 (N401, N389, N83, N177);
and AND4 (N402, N394, N397, N173, N221);
or OR3 (N403, N402, N281, N244);
not NOT1 (N404, N110);
nand NAND4 (N405, N393, N153, N164, N240);
and AND4 (N406, N405, N324, N230, N241);
xor XOR2 (N407, N400, N245);
or OR2 (N408, N399, N5);
buf BUF1 (N409, N407);
and AND3 (N410, N408, N32, N296);
and AND2 (N411, N406, N97);
and AND2 (N412, N392, N307);
or OR2 (N413, N403, N317);
and AND2 (N414, N395, N161);
not NOT1 (N415, N413);
or OR4 (N416, N409, N190, N153, N135);
nand NAND3 (N417, N396, N153, N385);
buf BUF1 (N418, N88);
xor XOR2 (N419, N404, N97);
buf BUF1 (N420, N415);
or OR3 (N421, N416, N29, N38);
xor XOR2 (N422, N418, N299);
nand NAND2 (N423, N401, N152);
not NOT1 (N424, N412);
nor NOR2 (N425, N422, N85);
xor XOR2 (N426, N411, N45);
not NOT1 (N427, N414);
and AND2 (N428, N421, N149);
xor XOR2 (N429, N410, N426);
xor XOR2 (N430, N72, N415);
or OR3 (N431, N423, N100, N206);
nand NAND2 (N432, N427, N212);
or OR2 (N433, N425, N23);
nor NOR2 (N434, N431, N113);
or OR2 (N435, N424, N208);
and AND4 (N436, N434, N237, N174, N310);
nand NAND3 (N437, N420, N149, N177);
nor NOR4 (N438, N436, N280, N106, N180);
and AND3 (N439, N433, N205, N364);
nor NOR3 (N440, N429, N239, N158);
and AND4 (N441, N435, N8, N418, N397);
nand NAND3 (N442, N437, N73, N174);
nor NOR2 (N443, N441, N114);
buf BUF1 (N444, N428);
nand NAND2 (N445, N419, N286);
and AND4 (N446, N417, N112, N58, N86);
buf BUF1 (N447, N440);
xor XOR2 (N448, N439, N331);
nor NOR2 (N449, N444, N157);
not NOT1 (N450, N448);
nor NOR2 (N451, N450, N253);
and AND3 (N452, N445, N337, N434);
and AND3 (N453, N446, N238, N12);
xor XOR2 (N454, N447, N251);
not NOT1 (N455, N453);
and AND4 (N456, N449, N144, N212, N167);
and AND2 (N457, N454, N100);
and AND4 (N458, N457, N201, N196, N445);
buf BUF1 (N459, N438);
buf BUF1 (N460, N458);
not NOT1 (N461, N460);
and AND4 (N462, N461, N197, N428, N394);
not NOT1 (N463, N459);
nor NOR4 (N464, N452, N267, N258, N69);
or OR4 (N465, N456, N405, N312, N165);
buf BUF1 (N466, N443);
nor NOR3 (N467, N451, N2, N43);
or OR2 (N468, N455, N184);
or OR3 (N469, N432, N114, N46);
buf BUF1 (N470, N467);
nor NOR4 (N471, N462, N149, N216, N407);
nor NOR4 (N472, N471, N449, N410, N90);
and AND4 (N473, N442, N363, N158, N219);
or OR4 (N474, N468, N352, N146, N236);
xor XOR2 (N475, N463, N177);
nand NAND2 (N476, N470, N434);
and AND2 (N477, N465, N420);
nor NOR3 (N478, N477, N191, N447);
nand NAND3 (N479, N472, N426, N132);
nand NAND3 (N480, N479, N432, N175);
not NOT1 (N481, N474);
nor NOR2 (N482, N466, N61);
buf BUF1 (N483, N469);
nor NOR4 (N484, N430, N423, N336, N294);
not NOT1 (N485, N481);
xor XOR2 (N486, N484, N279);
and AND2 (N487, N464, N193);
buf BUF1 (N488, N483);
xor XOR2 (N489, N480, N387);
not NOT1 (N490, N488);
nand NAND3 (N491, N482, N377, N7);
or OR2 (N492, N489, N263);
not NOT1 (N493, N486);
xor XOR2 (N494, N493, N210);
buf BUF1 (N495, N485);
xor XOR2 (N496, N476, N372);
nor NOR2 (N497, N496, N205);
and AND4 (N498, N494, N413, N60, N374);
nand NAND3 (N499, N498, N5, N119);
or OR4 (N500, N491, N35, N246, N291);
xor XOR2 (N501, N499, N234);
and AND3 (N502, N487, N387, N288);
buf BUF1 (N503, N495);
not NOT1 (N504, N502);
or OR2 (N505, N503, N471);
and AND4 (N506, N478, N164, N27, N281);
and AND3 (N507, N506, N402, N352);
and AND2 (N508, N473, N223);
not NOT1 (N509, N507);
or OR3 (N510, N504, N407, N499);
nand NAND4 (N511, N505, N452, N50, N371);
xor XOR2 (N512, N490, N20);
nor NOR4 (N513, N509, N505, N454, N54);
nor NOR3 (N514, N512, N333, N414);
xor XOR2 (N515, N511, N255);
or OR4 (N516, N501, N102, N214, N57);
and AND4 (N517, N516, N351, N128, N367);
or OR4 (N518, N500, N101, N50, N512);
not NOT1 (N519, N510);
or OR3 (N520, N518, N327, N63);
nand NAND4 (N521, N497, N475, N176, N124);
not NOT1 (N522, N35);
not NOT1 (N523, N521);
xor XOR2 (N524, N523, N511);
nand NAND2 (N525, N492, N44);
buf BUF1 (N526, N514);
xor XOR2 (N527, N508, N255);
nor NOR4 (N528, N517, N178, N304, N52);
or OR4 (N529, N528, N205, N241, N317);
and AND4 (N530, N513, N99, N489, N320);
or OR3 (N531, N519, N181, N213);
nand NAND4 (N532, N529, N488, N209, N338);
nand NAND4 (N533, N527, N25, N134, N475);
or OR4 (N534, N530, N225, N516, N342);
or OR2 (N535, N533, N449);
xor XOR2 (N536, N534, N150);
nand NAND2 (N537, N526, N458);
nor NOR3 (N538, N537, N361, N281);
or OR2 (N539, N525, N387);
not NOT1 (N540, N539);
or OR2 (N541, N522, N437);
xor XOR2 (N542, N515, N334);
nor NOR4 (N543, N531, N235, N115, N173);
and AND4 (N544, N541, N464, N497, N238);
nor NOR3 (N545, N542, N505, N153);
nand NAND2 (N546, N520, N161);
or OR3 (N547, N532, N176, N483);
xor XOR2 (N548, N524, N513);
buf BUF1 (N549, N535);
not NOT1 (N550, N549);
nor NOR4 (N551, N548, N113, N510, N450);
buf BUF1 (N552, N544);
and AND2 (N553, N536, N490);
buf BUF1 (N554, N552);
nand NAND2 (N555, N551, N146);
and AND3 (N556, N546, N272, N209);
xor XOR2 (N557, N554, N27);
nand NAND4 (N558, N556, N259, N276, N484);
nand NAND3 (N559, N543, N71, N505);
or OR4 (N560, N558, N34, N410, N396);
not NOT1 (N561, N540);
nor NOR2 (N562, N560, N487);
xor XOR2 (N563, N561, N455);
buf BUF1 (N564, N559);
buf BUF1 (N565, N564);
or OR2 (N566, N545, N549);
and AND4 (N567, N555, N93, N48, N253);
and AND3 (N568, N553, N464, N49);
or OR4 (N569, N538, N530, N307, N333);
buf BUF1 (N570, N562);
nand NAND2 (N571, N567, N294);
or OR2 (N572, N557, N148);
xor XOR2 (N573, N547, N527);
nor NOR2 (N574, N563, N549);
nand NAND2 (N575, N569, N179);
not NOT1 (N576, N550);
xor XOR2 (N577, N566, N385);
nand NAND2 (N578, N568, N341);
nor NOR3 (N579, N576, N11, N364);
nor NOR4 (N580, N578, N386, N185, N241);
or OR4 (N581, N572, N200, N238, N540);
buf BUF1 (N582, N571);
nor NOR3 (N583, N581, N256, N343);
nand NAND2 (N584, N579, N110);
or OR2 (N585, N573, N137);
nor NOR3 (N586, N585, N412, N34);
and AND2 (N587, N570, N330);
nand NAND2 (N588, N583, N125);
not NOT1 (N589, N565);
not NOT1 (N590, N580);
nand NAND2 (N591, N588, N463);
nand NAND4 (N592, N590, N366, N2, N561);
nand NAND3 (N593, N586, N527, N457);
xor XOR2 (N594, N587, N204);
or OR2 (N595, N577, N501);
buf BUF1 (N596, N592);
xor XOR2 (N597, N575, N569);
nor NOR2 (N598, N574, N349);
nor NOR4 (N599, N591, N77, N566, N508);
or OR4 (N600, N593, N335, N359, N505);
or OR4 (N601, N582, N480, N372, N143);
buf BUF1 (N602, N589);
nor NOR4 (N603, N599, N301, N344, N167);
buf BUF1 (N604, N594);
nor NOR4 (N605, N598, N177, N329, N214);
nor NOR4 (N606, N596, N93, N564, N280);
xor XOR2 (N607, N604, N475);
and AND3 (N608, N601, N587, N571);
or OR4 (N609, N595, N601, N158, N247);
xor XOR2 (N610, N603, N356);
buf BUF1 (N611, N584);
nor NOR4 (N612, N611, N155, N597, N446);
or OR3 (N613, N70, N563, N450);
nand NAND3 (N614, N605, N189, N455);
xor XOR2 (N615, N610, N102);
xor XOR2 (N616, N612, N172);
or OR3 (N617, N602, N246, N558);
buf BUF1 (N618, N613);
nor NOR3 (N619, N615, N127, N216);
xor XOR2 (N620, N616, N296);
xor XOR2 (N621, N617, N413);
nand NAND2 (N622, N619, N140);
buf BUF1 (N623, N606);
and AND4 (N624, N623, N457, N41, N283);
not NOT1 (N625, N607);
xor XOR2 (N626, N625, N181);
xor XOR2 (N627, N620, N405);
nor NOR2 (N628, N621, N111);
xor XOR2 (N629, N614, N346);
nand NAND4 (N630, N600, N332, N351, N207);
buf BUF1 (N631, N627);
nor NOR2 (N632, N631, N133);
xor XOR2 (N633, N608, N211);
and AND3 (N634, N632, N354, N491);
xor XOR2 (N635, N624, N141);
xor XOR2 (N636, N634, N10);
nor NOR4 (N637, N626, N479, N539, N118);
not NOT1 (N638, N609);
xor XOR2 (N639, N629, N611);
or OR3 (N640, N635, N323, N129);
and AND2 (N641, N636, N76);
buf BUF1 (N642, N633);
nor NOR3 (N643, N642, N607, N214);
buf BUF1 (N644, N630);
or OR2 (N645, N638, N325);
xor XOR2 (N646, N618, N581);
nor NOR3 (N647, N646, N65, N421);
buf BUF1 (N648, N637);
or OR2 (N649, N641, N93);
not NOT1 (N650, N644);
nor NOR4 (N651, N643, N395, N182, N348);
nand NAND2 (N652, N648, N112);
and AND2 (N653, N649, N195);
and AND4 (N654, N622, N206, N38, N424);
or OR3 (N655, N654, N545, N150);
nand NAND2 (N656, N628, N232);
nor NOR4 (N657, N653, N542, N125, N357);
xor XOR2 (N658, N647, N329);
buf BUF1 (N659, N658);
buf BUF1 (N660, N651);
nand NAND3 (N661, N659, N238, N292);
nor NOR2 (N662, N657, N46);
not NOT1 (N663, N656);
and AND2 (N664, N645, N447);
nor NOR2 (N665, N650, N207);
not NOT1 (N666, N661);
nor NOR2 (N667, N639, N544);
not NOT1 (N668, N664);
buf BUF1 (N669, N660);
nand NAND4 (N670, N667, N348, N659, N581);
or OR2 (N671, N662, N473);
buf BUF1 (N672, N671);
and AND3 (N673, N655, N49, N434);
nor NOR3 (N674, N669, N376, N563);
and AND2 (N675, N670, N511);
not NOT1 (N676, N674);
xor XOR2 (N677, N663, N46);
nor NOR4 (N678, N672, N243, N656, N370);
nand NAND2 (N679, N677, N652);
not NOT1 (N680, N181);
nand NAND4 (N681, N675, N230, N169, N300);
nor NOR2 (N682, N678, N404);
and AND3 (N683, N682, N321, N289);
or OR4 (N684, N673, N386, N1, N68);
nor NOR4 (N685, N681, N202, N325, N680);
or OR4 (N686, N420, N75, N275, N240);
or OR4 (N687, N640, N294, N74, N578);
buf BUF1 (N688, N683);
and AND3 (N689, N686, N407, N121);
nand NAND3 (N690, N688, N659, N423);
buf BUF1 (N691, N685);
not NOT1 (N692, N676);
nor NOR4 (N693, N687, N137, N35, N160);
not NOT1 (N694, N668);
buf BUF1 (N695, N684);
buf BUF1 (N696, N695);
not NOT1 (N697, N689);
nor NOR2 (N698, N697, N139);
xor XOR2 (N699, N694, N99);
not NOT1 (N700, N690);
buf BUF1 (N701, N679);
buf BUF1 (N702, N665);
xor XOR2 (N703, N699, N674);
xor XOR2 (N704, N691, N660);
and AND3 (N705, N698, N642, N447);
nand NAND4 (N706, N666, N104, N387, N156);
xor XOR2 (N707, N696, N436);
xor XOR2 (N708, N692, N550);
xor XOR2 (N709, N705, N37);
or OR2 (N710, N709, N166);
nor NOR4 (N711, N693, N165, N280, N364);
nor NOR3 (N712, N703, N564, N499);
buf BUF1 (N713, N712);
nor NOR4 (N714, N708, N497, N464, N415);
and AND2 (N715, N711, N156);
not NOT1 (N716, N715);
nor NOR2 (N717, N706, N462);
xor XOR2 (N718, N716, N102);
nor NOR4 (N719, N707, N476, N174, N2);
nand NAND2 (N720, N710, N198);
and AND4 (N721, N701, N334, N142, N65);
or OR2 (N722, N702, N384);
nand NAND4 (N723, N704, N21, N209, N167);
nor NOR2 (N724, N722, N355);
or OR4 (N725, N721, N343, N353, N692);
buf BUF1 (N726, N700);
or OR2 (N727, N717, N289);
and AND3 (N728, N727, N653, N189);
not NOT1 (N729, N725);
buf BUF1 (N730, N714);
xor XOR2 (N731, N728, N408);
nor NOR4 (N732, N718, N243, N245, N299);
buf BUF1 (N733, N732);
not NOT1 (N734, N726);
buf BUF1 (N735, N723);
xor XOR2 (N736, N730, N105);
buf BUF1 (N737, N733);
or OR2 (N738, N735, N47);
nor NOR2 (N739, N720, N725);
not NOT1 (N740, N738);
nor NOR3 (N741, N729, N608, N611);
and AND4 (N742, N741, N201, N419, N619);
xor XOR2 (N743, N736, N488);
buf BUF1 (N744, N731);
and AND2 (N745, N734, N531);
or OR3 (N746, N719, N523, N195);
not NOT1 (N747, N743);
not NOT1 (N748, N739);
nand NAND4 (N749, N747, N456, N723, N707);
and AND3 (N750, N737, N162, N199);
and AND4 (N751, N713, N8, N193, N600);
not NOT1 (N752, N749);
and AND2 (N753, N745, N485);
or OR3 (N754, N748, N135, N35);
not NOT1 (N755, N750);
not NOT1 (N756, N724);
or OR4 (N757, N744, N38, N197, N364);
nand NAND4 (N758, N742, N460, N363, N615);
nand NAND2 (N759, N746, N659);
nand NAND3 (N760, N740, N102, N70);
and AND2 (N761, N753, N482);
xor XOR2 (N762, N754, N245);
xor XOR2 (N763, N751, N297);
nand NAND3 (N764, N757, N505, N626);
buf BUF1 (N765, N760);
nor NOR3 (N766, N756, N644, N296);
and AND2 (N767, N765, N452);
xor XOR2 (N768, N762, N583);
xor XOR2 (N769, N766, N504);
or OR3 (N770, N759, N330, N532);
or OR3 (N771, N768, N427, N679);
nand NAND3 (N772, N755, N30, N704);
not NOT1 (N773, N763);
nor NOR2 (N774, N770, N118);
and AND2 (N775, N773, N672);
buf BUF1 (N776, N767);
xor XOR2 (N777, N772, N33);
or OR2 (N778, N758, N174);
or OR4 (N779, N764, N470, N750, N307);
or OR4 (N780, N776, N574, N715, N501);
not NOT1 (N781, N761);
not NOT1 (N782, N771);
buf BUF1 (N783, N774);
or OR2 (N784, N777, N738);
not NOT1 (N785, N752);
nor NOR3 (N786, N778, N104, N575);
or OR3 (N787, N769, N535, N220);
buf BUF1 (N788, N775);
or OR2 (N789, N787, N204);
buf BUF1 (N790, N784);
xor XOR2 (N791, N782, N592);
nor NOR2 (N792, N783, N718);
not NOT1 (N793, N789);
and AND4 (N794, N780, N738, N265, N260);
and AND3 (N795, N792, N352, N522);
buf BUF1 (N796, N790);
not NOT1 (N797, N786);
nand NAND4 (N798, N788, N336, N173, N543);
nor NOR3 (N799, N781, N478, N76);
and AND2 (N800, N797, N292);
not NOT1 (N801, N799);
xor XOR2 (N802, N801, N449);
and AND4 (N803, N794, N744, N793, N300);
buf BUF1 (N804, N254);
nand NAND2 (N805, N800, N733);
buf BUF1 (N806, N798);
or OR4 (N807, N802, N670, N706, N692);
xor XOR2 (N808, N795, N99);
buf BUF1 (N809, N806);
and AND4 (N810, N803, N95, N796, N278);
or OR2 (N811, N190, N533);
nor NOR3 (N812, N808, N26, N412);
or OR2 (N813, N804, N598);
and AND3 (N814, N779, N531, N717);
nand NAND3 (N815, N812, N50, N130);
buf BUF1 (N816, N791);
and AND3 (N817, N807, N511, N570);
buf BUF1 (N818, N785);
and AND4 (N819, N809, N52, N718, N599);
xor XOR2 (N820, N810, N192);
buf BUF1 (N821, N811);
xor XOR2 (N822, N813, N344);
and AND4 (N823, N822, N329, N811, N691);
nand NAND3 (N824, N815, N296, N705);
or OR3 (N825, N824, N497, N791);
or OR2 (N826, N817, N657);
or OR3 (N827, N818, N142, N340);
buf BUF1 (N828, N825);
xor XOR2 (N829, N819, N242);
and AND2 (N830, N828, N698);
or OR2 (N831, N829, N593);
buf BUF1 (N832, N823);
nand NAND2 (N833, N814, N360);
not NOT1 (N834, N833);
and AND3 (N835, N830, N269, N180);
or OR2 (N836, N821, N388);
nor NOR2 (N837, N836, N44);
and AND3 (N838, N834, N308, N142);
xor XOR2 (N839, N831, N673);
xor XOR2 (N840, N832, N688);
nor NOR3 (N841, N820, N416, N804);
not NOT1 (N842, N839);
or OR3 (N843, N840, N696, N143);
xor XOR2 (N844, N805, N624);
nand NAND3 (N845, N841, N108, N399);
and AND4 (N846, N835, N755, N479, N38);
and AND2 (N847, N826, N285);
nand NAND4 (N848, N844, N173, N595, N237);
nor NOR4 (N849, N838, N352, N670, N523);
nor NOR3 (N850, N827, N238, N33);
not NOT1 (N851, N816);
xor XOR2 (N852, N848, N314);
xor XOR2 (N853, N847, N591);
not NOT1 (N854, N852);
nor NOR3 (N855, N837, N717, N648);
or OR2 (N856, N846, N828);
buf BUF1 (N857, N842);
nor NOR2 (N858, N845, N825);
nand NAND4 (N859, N858, N411, N236, N692);
nand NAND3 (N860, N849, N822, N440);
or OR3 (N861, N854, N352, N497);
xor XOR2 (N862, N853, N323);
xor XOR2 (N863, N843, N317);
not NOT1 (N864, N861);
buf BUF1 (N865, N864);
xor XOR2 (N866, N862, N73);
not NOT1 (N867, N866);
or OR2 (N868, N867, N240);
or OR3 (N869, N868, N151, N795);
nor NOR4 (N870, N856, N70, N710, N815);
or OR3 (N871, N850, N620, N362);
and AND4 (N872, N859, N784, N466, N551);
nand NAND4 (N873, N872, N738, N761, N236);
nor NOR2 (N874, N871, N779);
or OR2 (N875, N870, N268);
buf BUF1 (N876, N855);
and AND2 (N877, N860, N628);
buf BUF1 (N878, N857);
nor NOR3 (N879, N877, N769, N203);
or OR2 (N880, N863, N59);
nor NOR4 (N881, N851, N690, N27, N259);
xor XOR2 (N882, N881, N283);
buf BUF1 (N883, N873);
or OR2 (N884, N865, N90);
and AND4 (N885, N869, N784, N331, N277);
nand NAND4 (N886, N884, N609, N413, N538);
xor XOR2 (N887, N875, N438);
not NOT1 (N888, N882);
and AND3 (N889, N880, N831, N827);
xor XOR2 (N890, N879, N749);
or OR3 (N891, N888, N538, N750);
nor NOR3 (N892, N890, N448, N583);
and AND2 (N893, N885, N872);
or OR2 (N894, N874, N484);
or OR3 (N895, N892, N231, N496);
not NOT1 (N896, N893);
buf BUF1 (N897, N896);
or OR4 (N898, N883, N154, N817, N373);
and AND4 (N899, N898, N809, N762, N96);
or OR4 (N900, N878, N466, N590, N452);
and AND3 (N901, N899, N821, N628);
nor NOR3 (N902, N901, N856, N684);
buf BUF1 (N903, N889);
nand NAND3 (N904, N887, N264, N794);
or OR2 (N905, N897, N569);
or OR2 (N906, N876, N40);
nand NAND3 (N907, N894, N228, N856);
nand NAND2 (N908, N904, N889);
nor NOR2 (N909, N907, N838);
nand NAND2 (N910, N908, N875);
nor NOR2 (N911, N910, N414);
or OR2 (N912, N891, N753);
or OR3 (N913, N903, N855, N400);
and AND2 (N914, N900, N757);
nor NOR3 (N915, N909, N310, N55);
nand NAND4 (N916, N886, N870, N358, N56);
not NOT1 (N917, N912);
not NOT1 (N918, N916);
and AND3 (N919, N914, N610, N572);
nand NAND3 (N920, N919, N291, N859);
buf BUF1 (N921, N905);
or OR2 (N922, N906, N411);
and AND3 (N923, N915, N717, N90);
xor XOR2 (N924, N918, N541);
xor XOR2 (N925, N920, N203);
nor NOR4 (N926, N913, N150, N305, N806);
not NOT1 (N927, N922);
xor XOR2 (N928, N923, N57);
or OR4 (N929, N911, N76, N526, N746);
nand NAND2 (N930, N927, N16);
or OR3 (N931, N924, N551, N849);
not NOT1 (N932, N902);
buf BUF1 (N933, N925);
nand NAND4 (N934, N930, N381, N700, N600);
or OR2 (N935, N928, N562);
nor NOR3 (N936, N932, N370, N129);
nand NAND4 (N937, N917, N164, N65, N622);
not NOT1 (N938, N937);
nand NAND2 (N939, N926, N211);
and AND2 (N940, N934, N45);
nor NOR2 (N941, N936, N913);
nand NAND4 (N942, N929, N566, N240, N477);
buf BUF1 (N943, N921);
xor XOR2 (N944, N940, N373);
and AND4 (N945, N941, N817, N944, N944);
nand NAND4 (N946, N676, N220, N568, N123);
buf BUF1 (N947, N931);
buf BUF1 (N948, N935);
or OR4 (N949, N939, N735, N63, N226);
nand NAND3 (N950, N895, N731, N683);
nand NAND3 (N951, N948, N253, N766);
buf BUF1 (N952, N938);
or OR3 (N953, N951, N425, N588);
not NOT1 (N954, N942);
and AND2 (N955, N945, N107);
buf BUF1 (N956, N953);
nor NOR3 (N957, N955, N661, N708);
not NOT1 (N958, N952);
not NOT1 (N959, N933);
xor XOR2 (N960, N949, N350);
or OR3 (N961, N956, N655, N637);
xor XOR2 (N962, N957, N697);
xor XOR2 (N963, N961, N772);
buf BUF1 (N964, N958);
nor NOR3 (N965, N954, N2, N318);
nor NOR4 (N966, N962, N302, N861, N450);
buf BUF1 (N967, N964);
buf BUF1 (N968, N946);
not NOT1 (N969, N963);
or OR2 (N970, N947, N317);
not NOT1 (N971, N943);
nor NOR2 (N972, N968, N71);
buf BUF1 (N973, N959);
nor NOR3 (N974, N971, N545, N661);
buf BUF1 (N975, N950);
xor XOR2 (N976, N975, N736);
nor NOR3 (N977, N976, N447, N521);
nor NOR2 (N978, N967, N597);
not NOT1 (N979, N974);
and AND3 (N980, N970, N973, N267);
not NOT1 (N981, N349);
buf BUF1 (N982, N981);
buf BUF1 (N983, N980);
nand NAND2 (N984, N966, N111);
nand NAND4 (N985, N984, N603, N355, N771);
xor XOR2 (N986, N972, N715);
not NOT1 (N987, N985);
or OR4 (N988, N969, N85, N884, N209);
xor XOR2 (N989, N982, N70);
xor XOR2 (N990, N977, N921);
and AND2 (N991, N965, N728);
xor XOR2 (N992, N979, N844);
or OR4 (N993, N983, N839, N741, N707);
nand NAND2 (N994, N988, N426);
or OR2 (N995, N960, N86);
not NOT1 (N996, N993);
or OR4 (N997, N986, N745, N633, N57);
or OR2 (N998, N978, N297);
and AND3 (N999, N996, N455, N407);
nor NOR3 (N1000, N995, N976, N105);
or OR2 (N1001, N998, N64);
or OR3 (N1002, N997, N282, N704);
xor XOR2 (N1003, N1001, N928);
nor NOR3 (N1004, N987, N831, N433);
nand NAND4 (N1005, N1000, N837, N155, N87);
nand NAND3 (N1006, N989, N232, N71);
or OR3 (N1007, N1002, N824, N154);
nor NOR4 (N1008, N994, N869, N577, N650);
nor NOR2 (N1009, N1003, N720);
nor NOR4 (N1010, N1005, N456, N605, N393);
and AND2 (N1011, N992, N101);
not NOT1 (N1012, N1004);
or OR2 (N1013, N991, N529);
nand NAND2 (N1014, N1006, N877);
nand NAND4 (N1015, N1011, N151, N37, N238);
nand NAND2 (N1016, N999, N655);
buf BUF1 (N1017, N1013);
nor NOR3 (N1018, N990, N499, N90);
or OR4 (N1019, N1007, N193, N233, N827);
or OR4 (N1020, N1014, N785, N610, N286);
not NOT1 (N1021, N1017);
nor NOR3 (N1022, N1018, N416, N829);
nand NAND3 (N1023, N1008, N482, N465);
xor XOR2 (N1024, N1022, N919);
and AND3 (N1025, N1015, N517, N940);
and AND4 (N1026, N1016, N131, N170, N48);
buf BUF1 (N1027, N1019);
nor NOR2 (N1028, N1023, N395);
nor NOR2 (N1029, N1009, N987);
not NOT1 (N1030, N1027);
nand NAND4 (N1031, N1020, N533, N132, N124);
or OR2 (N1032, N1031, N1028);
nor NOR4 (N1033, N814, N955, N679, N744);
buf BUF1 (N1034, N1025);
or OR4 (N1035, N1029, N565, N684, N739);
not NOT1 (N1036, N1035);
not NOT1 (N1037, N1034);
nor NOR4 (N1038, N1024, N787, N316, N1003);
and AND3 (N1039, N1037, N354, N1010);
or OR4 (N1040, N338, N203, N518, N173);
xor XOR2 (N1041, N1033, N502);
and AND4 (N1042, N1038, N794, N495, N591);
not NOT1 (N1043, N1012);
and AND2 (N1044, N1036, N285);
xor XOR2 (N1045, N1026, N833);
not NOT1 (N1046, N1030);
or OR3 (N1047, N1021, N989, N214);
not NOT1 (N1048, N1032);
nand NAND4 (N1049, N1042, N114, N336, N997);
buf BUF1 (N1050, N1044);
nor NOR3 (N1051, N1049, N383, N311);
or OR3 (N1052, N1043, N994, N915);
nor NOR3 (N1053, N1052, N661, N37);
nand NAND3 (N1054, N1047, N107, N276);
and AND4 (N1055, N1050, N908, N625, N202);
xor XOR2 (N1056, N1053, N803);
xor XOR2 (N1057, N1045, N1034);
or OR3 (N1058, N1041, N339, N370);
not NOT1 (N1059, N1056);
nor NOR2 (N1060, N1040, N634);
xor XOR2 (N1061, N1039, N37);
or OR2 (N1062, N1061, N649);
not NOT1 (N1063, N1062);
xor XOR2 (N1064, N1060, N108);
not NOT1 (N1065, N1059);
or OR4 (N1066, N1046, N452, N719, N960);
not NOT1 (N1067, N1065);
buf BUF1 (N1068, N1067);
buf BUF1 (N1069, N1066);
xor XOR2 (N1070, N1058, N852);
buf BUF1 (N1071, N1051);
or OR4 (N1072, N1048, N32, N141, N734);
and AND3 (N1073, N1055, N329, N37);
and AND3 (N1074, N1069, N416, N137);
xor XOR2 (N1075, N1064, N384);
or OR4 (N1076, N1054, N191, N415, N877);
nand NAND3 (N1077, N1073, N452, N995);
nor NOR4 (N1078, N1076, N274, N206, N792);
not NOT1 (N1079, N1068);
and AND4 (N1080, N1063, N546, N612, N387);
or OR4 (N1081, N1074, N1069, N28, N175);
not NOT1 (N1082, N1081);
xor XOR2 (N1083, N1077, N349);
xor XOR2 (N1084, N1070, N61);
not NOT1 (N1085, N1071);
not NOT1 (N1086, N1057);
or OR2 (N1087, N1086, N122);
xor XOR2 (N1088, N1072, N218);
xor XOR2 (N1089, N1075, N173);
or OR3 (N1090, N1083, N168, N651);
nor NOR4 (N1091, N1080, N793, N761, N909);
buf BUF1 (N1092, N1091);
nor NOR3 (N1093, N1090, N912, N307);
and AND2 (N1094, N1089, N477);
and AND4 (N1095, N1085, N320, N796, N1064);
buf BUF1 (N1096, N1084);
xor XOR2 (N1097, N1088, N598);
xor XOR2 (N1098, N1079, N1045);
nor NOR4 (N1099, N1096, N564, N283, N793);
nor NOR2 (N1100, N1082, N62);
nand NAND4 (N1101, N1087, N182, N942, N271);
nor NOR4 (N1102, N1078, N368, N631, N836);
and AND3 (N1103, N1101, N300, N917);
nand NAND3 (N1104, N1103, N406, N467);
nor NOR3 (N1105, N1102, N270, N1012);
nand NAND2 (N1106, N1098, N680);
or OR3 (N1107, N1097, N831, N308);
and AND3 (N1108, N1092, N215, N696);
nor NOR4 (N1109, N1105, N224, N858, N144);
not NOT1 (N1110, N1109);
buf BUF1 (N1111, N1099);
nand NAND2 (N1112, N1094, N198);
buf BUF1 (N1113, N1095);
nand NAND2 (N1114, N1100, N419);
not NOT1 (N1115, N1111);
and AND4 (N1116, N1093, N98, N225, N129);
buf BUF1 (N1117, N1108);
and AND3 (N1118, N1114, N940, N440);
and AND4 (N1119, N1106, N1105, N832, N955);
not NOT1 (N1120, N1113);
and AND2 (N1121, N1115, N766);
xor XOR2 (N1122, N1119, N502);
nand NAND3 (N1123, N1112, N1114, N842);
and AND3 (N1124, N1104, N392, N559);
xor XOR2 (N1125, N1121, N1014);
buf BUF1 (N1126, N1110);
buf BUF1 (N1127, N1122);
not NOT1 (N1128, N1127);
not NOT1 (N1129, N1125);
nor NOR2 (N1130, N1129, N281);
or OR4 (N1131, N1123, N855, N457, N86);
or OR2 (N1132, N1116, N264);
xor XOR2 (N1133, N1117, N208);
xor XOR2 (N1134, N1124, N986);
and AND4 (N1135, N1130, N208, N187, N91);
and AND4 (N1136, N1134, N591, N670, N958);
nand NAND3 (N1137, N1107, N45, N899);
or OR3 (N1138, N1128, N613, N350);
buf BUF1 (N1139, N1120);
nor NOR4 (N1140, N1137, N1117, N431, N37);
and AND3 (N1141, N1133, N975, N408);
not NOT1 (N1142, N1139);
nor NOR2 (N1143, N1118, N831);
not NOT1 (N1144, N1140);
xor XOR2 (N1145, N1144, N732);
or OR4 (N1146, N1138, N610, N52, N797);
or OR2 (N1147, N1141, N318);
nand NAND2 (N1148, N1146, N866);
nand NAND4 (N1149, N1132, N599, N513, N992);
and AND4 (N1150, N1126, N733, N446, N1034);
buf BUF1 (N1151, N1135);
nand NAND2 (N1152, N1136, N636);
and AND4 (N1153, N1149, N252, N853, N655);
nand NAND4 (N1154, N1153, N384, N155, N344);
xor XOR2 (N1155, N1143, N442);
nor NOR3 (N1156, N1147, N115, N153);
nor NOR2 (N1157, N1142, N910);
and AND2 (N1158, N1157, N785);
and AND2 (N1159, N1154, N922);
nand NAND3 (N1160, N1156, N377, N910);
buf BUF1 (N1161, N1158);
not NOT1 (N1162, N1148);
and AND2 (N1163, N1155, N146);
buf BUF1 (N1164, N1152);
not NOT1 (N1165, N1160);
not NOT1 (N1166, N1165);
buf BUF1 (N1167, N1151);
xor XOR2 (N1168, N1166, N780);
not NOT1 (N1169, N1131);
buf BUF1 (N1170, N1150);
nor NOR3 (N1171, N1164, N686, N893);
or OR2 (N1172, N1145, N455);
or OR3 (N1173, N1170, N381, N936);
not NOT1 (N1174, N1169);
nor NOR2 (N1175, N1162, N700);
not NOT1 (N1176, N1174);
nor NOR4 (N1177, N1172, N1082, N970, N913);
xor XOR2 (N1178, N1167, N100);
xor XOR2 (N1179, N1159, N474);
not NOT1 (N1180, N1179);
nor NOR2 (N1181, N1163, N776);
buf BUF1 (N1182, N1175);
and AND3 (N1183, N1177, N686, N376);
xor XOR2 (N1184, N1168, N1026);
nor NOR3 (N1185, N1184, N437, N777);
not NOT1 (N1186, N1180);
or OR2 (N1187, N1176, N529);
xor XOR2 (N1188, N1173, N1138);
not NOT1 (N1189, N1183);
nand NAND4 (N1190, N1189, N195, N498, N1017);
buf BUF1 (N1191, N1181);
or OR4 (N1192, N1191, N383, N1134, N733);
buf BUF1 (N1193, N1192);
and AND3 (N1194, N1178, N162, N195);
and AND4 (N1195, N1186, N957, N1117, N329);
xor XOR2 (N1196, N1194, N816);
and AND2 (N1197, N1190, N970);
nor NOR3 (N1198, N1187, N30, N295);
xor XOR2 (N1199, N1193, N475);
nand NAND2 (N1200, N1161, N85);
or OR3 (N1201, N1199, N1000, N1149);
or OR4 (N1202, N1198, N992, N75, N910);
nand NAND4 (N1203, N1196, N169, N953, N974);
nor NOR4 (N1204, N1202, N937, N208, N200);
or OR4 (N1205, N1203, N209, N521, N854);
not NOT1 (N1206, N1171);
nand NAND4 (N1207, N1185, N598, N343, N1097);
nor NOR2 (N1208, N1195, N1073);
nor NOR2 (N1209, N1204, N606);
xor XOR2 (N1210, N1207, N622);
not NOT1 (N1211, N1201);
nor NOR2 (N1212, N1208, N597);
and AND2 (N1213, N1206, N953);
and AND2 (N1214, N1209, N579);
not NOT1 (N1215, N1205);
buf BUF1 (N1216, N1200);
and AND4 (N1217, N1216, N939, N348, N313);
buf BUF1 (N1218, N1212);
or OR3 (N1219, N1215, N865, N932);
and AND3 (N1220, N1217, N534, N346);
or OR3 (N1221, N1213, N993, N743);
nand NAND2 (N1222, N1214, N953);
nor NOR2 (N1223, N1220, N670);
buf BUF1 (N1224, N1211);
nor NOR4 (N1225, N1197, N1155, N985, N1050);
or OR2 (N1226, N1210, N1113);
xor XOR2 (N1227, N1219, N1095);
nand NAND3 (N1228, N1223, N727, N130);
buf BUF1 (N1229, N1218);
or OR2 (N1230, N1226, N376);
nor NOR4 (N1231, N1224, N215, N971, N1078);
xor XOR2 (N1232, N1230, N36);
xor XOR2 (N1233, N1225, N862);
not NOT1 (N1234, N1182);
and AND2 (N1235, N1232, N381);
nand NAND4 (N1236, N1228, N1133, N329, N1197);
nand NAND2 (N1237, N1188, N1021);
or OR2 (N1238, N1233, N638);
or OR2 (N1239, N1238, N199);
or OR4 (N1240, N1231, N620, N171, N980);
xor XOR2 (N1241, N1236, N188);
not NOT1 (N1242, N1235);
and AND3 (N1243, N1227, N588, N1031);
and AND3 (N1244, N1241, N696, N1115);
or OR2 (N1245, N1239, N641);
and AND2 (N1246, N1240, N1173);
nor NOR3 (N1247, N1221, N1146, N591);
nand NAND4 (N1248, N1246, N1122, N1062, N17);
or OR4 (N1249, N1242, N789, N726, N287);
not NOT1 (N1250, N1248);
buf BUF1 (N1251, N1247);
nand NAND4 (N1252, N1249, N71, N836, N22);
and AND4 (N1253, N1237, N745, N999, N566);
nand NAND3 (N1254, N1234, N364, N955);
xor XOR2 (N1255, N1222, N699);
and AND3 (N1256, N1253, N396, N823);
or OR3 (N1257, N1229, N794, N247);
not NOT1 (N1258, N1250);
not NOT1 (N1259, N1245);
nand NAND4 (N1260, N1244, N985, N541, N893);
nor NOR2 (N1261, N1243, N392);
or OR2 (N1262, N1255, N501);
and AND3 (N1263, N1261, N818, N344);
and AND4 (N1264, N1256, N1134, N1158, N220);
nor NOR3 (N1265, N1251, N790, N890);
not NOT1 (N1266, N1264);
not NOT1 (N1267, N1263);
nor NOR2 (N1268, N1259, N1072);
buf BUF1 (N1269, N1260);
xor XOR2 (N1270, N1269, N1143);
xor XOR2 (N1271, N1252, N588);
not NOT1 (N1272, N1271);
nor NOR2 (N1273, N1258, N236);
buf BUF1 (N1274, N1268);
nor NOR2 (N1275, N1257, N307);
buf BUF1 (N1276, N1265);
buf BUF1 (N1277, N1270);
or OR4 (N1278, N1262, N740, N475, N1213);
nand NAND3 (N1279, N1267, N160, N1230);
and AND3 (N1280, N1279, N816, N198);
not NOT1 (N1281, N1276);
and AND3 (N1282, N1254, N925, N963);
buf BUF1 (N1283, N1280);
not NOT1 (N1284, N1273);
or OR4 (N1285, N1284, N1146, N57, N1210);
not NOT1 (N1286, N1278);
nand NAND2 (N1287, N1277, N820);
or OR2 (N1288, N1285, N384);
nor NOR4 (N1289, N1282, N865, N817, N383);
and AND4 (N1290, N1281, N53, N710, N834);
nor NOR4 (N1291, N1289, N692, N698, N324);
buf BUF1 (N1292, N1288);
xor XOR2 (N1293, N1283, N617);
xor XOR2 (N1294, N1287, N584);
and AND3 (N1295, N1294, N601, N1083);
not NOT1 (N1296, N1293);
and AND3 (N1297, N1291, N701, N811);
nand NAND4 (N1298, N1297, N1121, N1045, N1188);
or OR3 (N1299, N1298, N908, N531);
nor NOR3 (N1300, N1295, N188, N1213);
nor NOR2 (N1301, N1299, N844);
nor NOR4 (N1302, N1274, N254, N437, N752);
nor NOR2 (N1303, N1286, N550);
xor XOR2 (N1304, N1275, N112);
buf BUF1 (N1305, N1303);
and AND4 (N1306, N1290, N496, N663, N1270);
not NOT1 (N1307, N1300);
nand NAND2 (N1308, N1296, N1272);
nor NOR4 (N1309, N934, N420, N73, N797);
buf BUF1 (N1310, N1266);
nor NOR3 (N1311, N1305, N451, N990);
buf BUF1 (N1312, N1301);
and AND3 (N1313, N1292, N558, N1231);
nand NAND2 (N1314, N1304, N610);
nor NOR3 (N1315, N1309, N8, N891);
and AND4 (N1316, N1310, N1310, N539, N1058);
nor NOR2 (N1317, N1316, N1103);
xor XOR2 (N1318, N1313, N819);
xor XOR2 (N1319, N1315, N307);
buf BUF1 (N1320, N1302);
or OR4 (N1321, N1320, N276, N981, N1023);
not NOT1 (N1322, N1307);
nor NOR3 (N1323, N1312, N664, N348);
not NOT1 (N1324, N1319);
nand NAND4 (N1325, N1318, N111, N1318, N154);
not NOT1 (N1326, N1317);
not NOT1 (N1327, N1326);
xor XOR2 (N1328, N1321, N1064);
and AND3 (N1329, N1308, N707, N1175);
nand NAND3 (N1330, N1324, N684, N410);
not NOT1 (N1331, N1311);
nor NOR2 (N1332, N1328, N1171);
nor NOR2 (N1333, N1322, N1160);
xor XOR2 (N1334, N1306, N1256);
buf BUF1 (N1335, N1333);
or OR2 (N1336, N1335, N1272);
not NOT1 (N1337, N1323);
buf BUF1 (N1338, N1331);
xor XOR2 (N1339, N1337, N433);
or OR4 (N1340, N1330, N1283, N1203, N796);
and AND2 (N1341, N1340, N573);
or OR2 (N1342, N1341, N1070);
xor XOR2 (N1343, N1342, N704);
buf BUF1 (N1344, N1329);
nand NAND3 (N1345, N1325, N684, N40);
xor XOR2 (N1346, N1336, N74);
and AND4 (N1347, N1338, N493, N1336, N843);
not NOT1 (N1348, N1332);
or OR3 (N1349, N1334, N835, N738);
nand NAND4 (N1350, N1327, N203, N695, N999);
buf BUF1 (N1351, N1314);
or OR3 (N1352, N1343, N159, N768);
and AND4 (N1353, N1351, N1031, N454, N386);
not NOT1 (N1354, N1352);
xor XOR2 (N1355, N1345, N49);
or OR3 (N1356, N1354, N156, N399);
buf BUF1 (N1357, N1350);
buf BUF1 (N1358, N1347);
or OR2 (N1359, N1353, N429);
buf BUF1 (N1360, N1355);
buf BUF1 (N1361, N1339);
nor NOR3 (N1362, N1344, N1023, N1117);
buf BUF1 (N1363, N1356);
or OR3 (N1364, N1358, N81, N822);
and AND4 (N1365, N1364, N986, N842, N163);
buf BUF1 (N1366, N1346);
and AND2 (N1367, N1360, N28);
nor NOR2 (N1368, N1349, N1127);
not NOT1 (N1369, N1365);
or OR3 (N1370, N1367, N318, N1208);
nand NAND4 (N1371, N1368, N212, N772, N850);
not NOT1 (N1372, N1371);
not NOT1 (N1373, N1357);
or OR3 (N1374, N1348, N475, N443);
not NOT1 (N1375, N1362);
not NOT1 (N1376, N1375);
nor NOR3 (N1377, N1361, N858, N333);
not NOT1 (N1378, N1363);
nand NAND2 (N1379, N1378, N1307);
nand NAND3 (N1380, N1359, N197, N1348);
nor NOR3 (N1381, N1369, N1234, N92);
or OR3 (N1382, N1366, N420, N1310);
xor XOR2 (N1383, N1373, N239);
nor NOR4 (N1384, N1370, N819, N293, N533);
nor NOR2 (N1385, N1382, N776);
buf BUF1 (N1386, N1384);
xor XOR2 (N1387, N1381, N603);
nor NOR4 (N1388, N1379, N1245, N112, N563);
xor XOR2 (N1389, N1372, N891);
buf BUF1 (N1390, N1380);
not NOT1 (N1391, N1390);
nor NOR4 (N1392, N1377, N1206, N438, N1000);
buf BUF1 (N1393, N1383);
nor NOR3 (N1394, N1376, N166, N461);
not NOT1 (N1395, N1386);
buf BUF1 (N1396, N1385);
nor NOR2 (N1397, N1392, N183);
or OR4 (N1398, N1397, N1023, N877, N789);
buf BUF1 (N1399, N1396);
nor NOR3 (N1400, N1374, N5, N244);
not NOT1 (N1401, N1389);
nor NOR4 (N1402, N1394, N203, N846, N454);
nor NOR2 (N1403, N1399, N1041);
xor XOR2 (N1404, N1403, N417);
nor NOR4 (N1405, N1401, N1221, N926, N683);
or OR2 (N1406, N1404, N95);
buf BUF1 (N1407, N1398);
not NOT1 (N1408, N1388);
or OR2 (N1409, N1387, N69);
and AND2 (N1410, N1400, N341);
not NOT1 (N1411, N1406);
buf BUF1 (N1412, N1391);
not NOT1 (N1413, N1402);
and AND3 (N1414, N1409, N1182, N151);
and AND2 (N1415, N1405, N393);
or OR4 (N1416, N1413, N786, N17, N680);
or OR3 (N1417, N1415, N1130, N584);
nand NAND3 (N1418, N1412, N667, N1015);
xor XOR2 (N1419, N1417, N789);
xor XOR2 (N1420, N1416, N530);
nor NOR3 (N1421, N1411, N640, N514);
nor NOR4 (N1422, N1395, N490, N465, N1067);
xor XOR2 (N1423, N1421, N1160);
buf BUF1 (N1424, N1408);
xor XOR2 (N1425, N1424, N1422);
and AND2 (N1426, N248, N1372);
not NOT1 (N1427, N1393);
nor NOR2 (N1428, N1418, N558);
nor NOR2 (N1429, N1427, N1020);
buf BUF1 (N1430, N1414);
not NOT1 (N1431, N1425);
nor NOR3 (N1432, N1410, N24, N1416);
nor NOR3 (N1433, N1426, N364, N319);
xor XOR2 (N1434, N1423, N1056);
and AND2 (N1435, N1434, N450);
xor XOR2 (N1436, N1435, N593);
nand NAND4 (N1437, N1429, N319, N997, N993);
nor NOR3 (N1438, N1437, N784, N1426);
not NOT1 (N1439, N1431);
buf BUF1 (N1440, N1419);
not NOT1 (N1441, N1407);
xor XOR2 (N1442, N1438, N760);
xor XOR2 (N1443, N1428, N1058);
not NOT1 (N1444, N1439);
nand NAND3 (N1445, N1441, N1164, N72);
not NOT1 (N1446, N1420);
and AND2 (N1447, N1432, N367);
not NOT1 (N1448, N1442);
or OR3 (N1449, N1445, N937, N161);
nor NOR4 (N1450, N1440, N124, N1167, N587);
nand NAND3 (N1451, N1436, N936, N1344);
xor XOR2 (N1452, N1448, N497);
not NOT1 (N1453, N1451);
nand NAND3 (N1454, N1450, N440, N6);
or OR3 (N1455, N1454, N383, N1327);
xor XOR2 (N1456, N1452, N111);
xor XOR2 (N1457, N1444, N1301);
xor XOR2 (N1458, N1430, N522);
xor XOR2 (N1459, N1433, N1361);
nor NOR3 (N1460, N1453, N1339, N860);
nand NAND4 (N1461, N1443, N1424, N858, N359);
or OR3 (N1462, N1449, N676, N549);
xor XOR2 (N1463, N1446, N151);
nor NOR4 (N1464, N1458, N1439, N1199, N3);
xor XOR2 (N1465, N1447, N1403);
or OR4 (N1466, N1459, N225, N1050, N376);
buf BUF1 (N1467, N1465);
xor XOR2 (N1468, N1460, N689);
nand NAND3 (N1469, N1467, N1254, N492);
nand NAND4 (N1470, N1468, N1194, N651, N536);
or OR2 (N1471, N1470, N1459);
not NOT1 (N1472, N1471);
nor NOR3 (N1473, N1472, N545, N502);
buf BUF1 (N1474, N1469);
not NOT1 (N1475, N1464);
and AND3 (N1476, N1462, N1376, N94);
xor XOR2 (N1477, N1466, N1185);
buf BUF1 (N1478, N1461);
or OR2 (N1479, N1463, N1390);
buf BUF1 (N1480, N1457);
xor XOR2 (N1481, N1473, N458);
xor XOR2 (N1482, N1478, N1144);
or OR4 (N1483, N1477, N436, N11, N1227);
nor NOR2 (N1484, N1455, N940);
or OR4 (N1485, N1476, N1269, N14, N913);
and AND4 (N1486, N1482, N1438, N823, N1314);
and AND4 (N1487, N1483, N1152, N632, N855);
and AND4 (N1488, N1485, N1396, N655, N974);
nor NOR2 (N1489, N1474, N855);
buf BUF1 (N1490, N1456);
xor XOR2 (N1491, N1484, N1160);
xor XOR2 (N1492, N1481, N846);
nor NOR4 (N1493, N1488, N314, N306, N511);
xor XOR2 (N1494, N1490, N882);
nand NAND2 (N1495, N1475, N738);
nand NAND4 (N1496, N1494, N747, N375, N237);
not NOT1 (N1497, N1492);
and AND4 (N1498, N1486, N743, N573, N864);
and AND2 (N1499, N1491, N308);
and AND4 (N1500, N1489, N44, N1001, N630);
not NOT1 (N1501, N1480);
or OR3 (N1502, N1499, N1374, N1204);
nor NOR2 (N1503, N1502, N1174);
nand NAND2 (N1504, N1479, N1503);
and AND4 (N1505, N887, N197, N765, N1432);
nand NAND2 (N1506, N1505, N931);
nand NAND3 (N1507, N1501, N371, N423);
and AND4 (N1508, N1498, N1485, N438, N1071);
not NOT1 (N1509, N1493);
and AND3 (N1510, N1497, N748, N1108);
or OR2 (N1511, N1509, N1468);
not NOT1 (N1512, N1500);
buf BUF1 (N1513, N1510);
and AND4 (N1514, N1508, N614, N55, N459);
buf BUF1 (N1515, N1506);
buf BUF1 (N1516, N1514);
not NOT1 (N1517, N1512);
xor XOR2 (N1518, N1487, N173);
nor NOR4 (N1519, N1513, N1193, N253, N1215);
nand NAND3 (N1520, N1507, N1314, N465);
xor XOR2 (N1521, N1511, N224);
not NOT1 (N1522, N1519);
not NOT1 (N1523, N1504);
nand NAND4 (N1524, N1495, N299, N1179, N978);
buf BUF1 (N1525, N1515);
buf BUF1 (N1526, N1525);
nand NAND2 (N1527, N1521, N460);
or OR2 (N1528, N1522, N627);
nand NAND2 (N1529, N1524, N167);
nand NAND4 (N1530, N1526, N1491, N1097, N166);
xor XOR2 (N1531, N1496, N716);
or OR2 (N1532, N1528, N218);
not NOT1 (N1533, N1531);
or OR4 (N1534, N1532, N686, N1251, N669);
or OR3 (N1535, N1517, N321, N563);
buf BUF1 (N1536, N1534);
and AND4 (N1537, N1536, N1059, N1508, N748);
nor NOR2 (N1538, N1530, N141);
and AND4 (N1539, N1529, N1510, N1301, N1020);
xor XOR2 (N1540, N1533, N500);
nor NOR2 (N1541, N1516, N837);
buf BUF1 (N1542, N1518);
nand NAND4 (N1543, N1539, N1182, N811, N129);
and AND4 (N1544, N1541, N1433, N388, N199);
and AND2 (N1545, N1542, N1291);
or OR3 (N1546, N1520, N537, N786);
nand NAND3 (N1547, N1540, N568, N474);
not NOT1 (N1548, N1538);
buf BUF1 (N1549, N1537);
nor NOR4 (N1550, N1535, N578, N1368, N353);
xor XOR2 (N1551, N1545, N1016);
nor NOR2 (N1552, N1548, N123);
buf BUF1 (N1553, N1544);
not NOT1 (N1554, N1550);
not NOT1 (N1555, N1553);
and AND3 (N1556, N1547, N1062, N607);
not NOT1 (N1557, N1556);
and AND2 (N1558, N1523, N103);
nand NAND4 (N1559, N1552, N48, N592, N1447);
and AND4 (N1560, N1558, N1297, N141, N690);
nor NOR3 (N1561, N1549, N1303, N726);
nor NOR3 (N1562, N1543, N48, N1260);
nand NAND2 (N1563, N1546, N746);
not NOT1 (N1564, N1557);
nand NAND2 (N1565, N1560, N1432);
not NOT1 (N1566, N1555);
buf BUF1 (N1567, N1561);
xor XOR2 (N1568, N1559, N1018);
not NOT1 (N1569, N1566);
nand NAND2 (N1570, N1564, N969);
nor NOR2 (N1571, N1551, N253);
buf BUF1 (N1572, N1567);
nand NAND2 (N1573, N1563, N789);
not NOT1 (N1574, N1570);
buf BUF1 (N1575, N1572);
xor XOR2 (N1576, N1574, N1521);
nor NOR4 (N1577, N1575, N810, N1305, N1183);
xor XOR2 (N1578, N1554, N785);
not NOT1 (N1579, N1569);
nand NAND4 (N1580, N1576, N815, N1572, N613);
nand NAND3 (N1581, N1562, N620, N739);
nand NAND4 (N1582, N1527, N1042, N483, N549);
xor XOR2 (N1583, N1571, N1031);
not NOT1 (N1584, N1580);
nand NAND2 (N1585, N1579, N1473);
nand NAND3 (N1586, N1568, N991, N643);
and AND2 (N1587, N1585, N987);
not NOT1 (N1588, N1583);
not NOT1 (N1589, N1577);
nor NOR4 (N1590, N1587, N712, N525, N1152);
nor NOR2 (N1591, N1586, N82);
xor XOR2 (N1592, N1584, N329);
xor XOR2 (N1593, N1589, N335);
nand NAND3 (N1594, N1590, N229, N601);
nand NAND2 (N1595, N1581, N637);
nor NOR3 (N1596, N1588, N389, N1283);
nor NOR2 (N1597, N1565, N675);
and AND4 (N1598, N1592, N1500, N768, N911);
nand NAND3 (N1599, N1595, N892, N1385);
xor XOR2 (N1600, N1591, N366);
nor NOR2 (N1601, N1598, N24);
and AND3 (N1602, N1573, N1202, N207);
or OR2 (N1603, N1600, N951);
or OR3 (N1604, N1601, N116, N270);
not NOT1 (N1605, N1604);
or OR4 (N1606, N1599, N1374, N133, N1230);
nand NAND2 (N1607, N1593, N839);
and AND4 (N1608, N1603, N1273, N1224, N444);
and AND4 (N1609, N1578, N1486, N1034, N896);
and AND4 (N1610, N1609, N1038, N298, N536);
not NOT1 (N1611, N1594);
not NOT1 (N1612, N1605);
and AND3 (N1613, N1606, N726, N1031);
xor XOR2 (N1614, N1611, N1295);
nand NAND3 (N1615, N1613, N82, N1332);
xor XOR2 (N1616, N1614, N1337);
xor XOR2 (N1617, N1597, N625);
nand NAND3 (N1618, N1607, N599, N318);
buf BUF1 (N1619, N1608);
not NOT1 (N1620, N1612);
not NOT1 (N1621, N1620);
xor XOR2 (N1622, N1618, N897);
buf BUF1 (N1623, N1617);
buf BUF1 (N1624, N1619);
xor XOR2 (N1625, N1602, N1222);
buf BUF1 (N1626, N1624);
xor XOR2 (N1627, N1610, N1473);
nor NOR4 (N1628, N1625, N261, N421, N258);
not NOT1 (N1629, N1628);
buf BUF1 (N1630, N1629);
or OR4 (N1631, N1622, N605, N305, N702);
and AND2 (N1632, N1621, N976);
not NOT1 (N1633, N1615);
nand NAND4 (N1634, N1626, N1096, N840, N646);
nor NOR2 (N1635, N1630, N287);
or OR3 (N1636, N1596, N1500, N841);
and AND2 (N1637, N1582, N854);
nand NAND3 (N1638, N1627, N518, N820);
or OR3 (N1639, N1634, N1364, N1295);
and AND4 (N1640, N1638, N11, N613, N1500);
nor NOR3 (N1641, N1635, N1212, N719);
nor NOR3 (N1642, N1640, N57, N602);
and AND4 (N1643, N1637, N1167, N965, N707);
or OR2 (N1644, N1641, N533);
and AND3 (N1645, N1632, N246, N931);
and AND4 (N1646, N1639, N1091, N1113, N796);
nor NOR4 (N1647, N1642, N100, N221, N1497);
and AND4 (N1648, N1647, N1535, N685, N1561);
and AND2 (N1649, N1633, N195);
buf BUF1 (N1650, N1623);
nand NAND2 (N1651, N1645, N1377);
or OR2 (N1652, N1643, N163);
or OR4 (N1653, N1648, N1399, N684, N1349);
not NOT1 (N1654, N1636);
or OR2 (N1655, N1649, N417);
xor XOR2 (N1656, N1616, N1207);
xor XOR2 (N1657, N1644, N1098);
or OR4 (N1658, N1651, N256, N1389, N722);
buf BUF1 (N1659, N1658);
buf BUF1 (N1660, N1657);
buf BUF1 (N1661, N1659);
and AND4 (N1662, N1631, N1385, N1552, N1631);
buf BUF1 (N1663, N1646);
buf BUF1 (N1664, N1653);
nor NOR4 (N1665, N1662, N1594, N173, N648);
nor NOR3 (N1666, N1660, N149, N1232);
xor XOR2 (N1667, N1661, N1331);
or OR3 (N1668, N1655, N915, N630);
buf BUF1 (N1669, N1652);
and AND4 (N1670, N1654, N626, N906, N1586);
and AND4 (N1671, N1665, N647, N289, N1385);
buf BUF1 (N1672, N1664);
or OR2 (N1673, N1650, N1308);
nor NOR2 (N1674, N1673, N1305);
or OR3 (N1675, N1667, N592, N157);
nand NAND4 (N1676, N1672, N786, N1262, N316);
nand NAND4 (N1677, N1656, N323, N718, N1111);
nor NOR4 (N1678, N1675, N229, N192, N387);
nand NAND2 (N1679, N1669, N523);
and AND4 (N1680, N1666, N399, N1406, N320);
xor XOR2 (N1681, N1663, N64);
buf BUF1 (N1682, N1681);
nand NAND3 (N1683, N1676, N34, N832);
not NOT1 (N1684, N1668);
or OR4 (N1685, N1679, N1122, N1319, N221);
or OR3 (N1686, N1685, N189, N312);
nand NAND4 (N1687, N1686, N639, N1646, N1217);
nand NAND3 (N1688, N1683, N888, N450);
xor XOR2 (N1689, N1684, N1192);
not NOT1 (N1690, N1674);
not NOT1 (N1691, N1687);
nor NOR4 (N1692, N1688, N1384, N304, N714);
nor NOR3 (N1693, N1671, N381, N1478);
and AND4 (N1694, N1689, N883, N267, N663);
nand NAND4 (N1695, N1678, N1691, N1196, N1325);
xor XOR2 (N1696, N1581, N578);
xor XOR2 (N1697, N1680, N805);
and AND3 (N1698, N1692, N1361, N1572);
xor XOR2 (N1699, N1690, N1375);
not NOT1 (N1700, N1693);
xor XOR2 (N1701, N1700, N545);
or OR2 (N1702, N1677, N895);
nor NOR2 (N1703, N1696, N1675);
or OR4 (N1704, N1703, N1569, N1378, N8);
nand NAND3 (N1705, N1697, N202, N1561);
xor XOR2 (N1706, N1694, N701);
or OR4 (N1707, N1670, N689, N673, N1005);
not NOT1 (N1708, N1705);
buf BUF1 (N1709, N1699);
nor NOR4 (N1710, N1695, N992, N854, N682);
and AND2 (N1711, N1682, N1374);
not NOT1 (N1712, N1707);
xor XOR2 (N1713, N1711, N1214);
or OR4 (N1714, N1712, N355, N292, N262);
nand NAND3 (N1715, N1706, N1539, N673);
not NOT1 (N1716, N1702);
buf BUF1 (N1717, N1716);
xor XOR2 (N1718, N1704, N595);
not NOT1 (N1719, N1710);
not NOT1 (N1720, N1714);
nor NOR4 (N1721, N1719, N916, N1715, N359);
not NOT1 (N1722, N878);
and AND2 (N1723, N1722, N1042);
buf BUF1 (N1724, N1698);
and AND2 (N1725, N1713, N28);
nor NOR3 (N1726, N1724, N806, N1193);
nor NOR2 (N1727, N1720, N579);
or OR3 (N1728, N1709, N926, N1110);
or OR3 (N1729, N1727, N87, N430);
nand NAND2 (N1730, N1723, N520);
buf BUF1 (N1731, N1701);
not NOT1 (N1732, N1717);
nor NOR2 (N1733, N1721, N644);
and AND3 (N1734, N1731, N127, N1592);
nor NOR2 (N1735, N1734, N82);
buf BUF1 (N1736, N1708);
xor XOR2 (N1737, N1728, N899);
nor NOR2 (N1738, N1737, N1510);
xor XOR2 (N1739, N1718, N1517);
xor XOR2 (N1740, N1739, N1612);
or OR3 (N1741, N1730, N575, N885);
xor XOR2 (N1742, N1726, N463);
nand NAND4 (N1743, N1738, N981, N979, N228);
and AND2 (N1744, N1729, N1011);
and AND4 (N1745, N1742, N697, N585, N325);
not NOT1 (N1746, N1736);
or OR3 (N1747, N1732, N79, N648);
not NOT1 (N1748, N1741);
or OR4 (N1749, N1746, N938, N102, N1327);
not NOT1 (N1750, N1725);
not NOT1 (N1751, N1733);
nor NOR2 (N1752, N1744, N448);
and AND3 (N1753, N1740, N1054, N477);
nor NOR4 (N1754, N1745, N1702, N929, N930);
and AND3 (N1755, N1735, N275, N630);
nand NAND4 (N1756, N1748, N770, N588, N860);
nor NOR3 (N1757, N1755, N229, N14);
buf BUF1 (N1758, N1743);
xor XOR2 (N1759, N1756, N1584);
nor NOR4 (N1760, N1752, N1562, N1177, N213);
and AND4 (N1761, N1750, N328, N774, N999);
nand NAND3 (N1762, N1757, N908, N1040);
nand NAND4 (N1763, N1754, N687, N917, N584);
xor XOR2 (N1764, N1761, N1462);
buf BUF1 (N1765, N1747);
not NOT1 (N1766, N1760);
not NOT1 (N1767, N1758);
nand NAND4 (N1768, N1766, N323, N1092, N1325);
nor NOR3 (N1769, N1751, N1686, N417);
and AND3 (N1770, N1767, N8, N467);
not NOT1 (N1771, N1749);
buf BUF1 (N1772, N1763);
nor NOR4 (N1773, N1759, N734, N1759, N1731);
or OR2 (N1774, N1764, N358);
or OR3 (N1775, N1753, N1319, N447);
nor NOR3 (N1776, N1772, N1258, N478);
nor NOR2 (N1777, N1765, N635);
nor NOR3 (N1778, N1768, N154, N809);
buf BUF1 (N1779, N1775);
buf BUF1 (N1780, N1773);
xor XOR2 (N1781, N1770, N1083);
or OR2 (N1782, N1779, N1647);
xor XOR2 (N1783, N1780, N903);
not NOT1 (N1784, N1771);
and AND2 (N1785, N1776, N158);
nor NOR3 (N1786, N1774, N744, N1443);
and AND2 (N1787, N1777, N1124);
nor NOR3 (N1788, N1782, N1528, N901);
xor XOR2 (N1789, N1783, N805);
not NOT1 (N1790, N1784);
nor NOR2 (N1791, N1762, N1479);
nor NOR4 (N1792, N1786, N51, N966, N1157);
and AND2 (N1793, N1785, N995);
nor NOR2 (N1794, N1793, N738);
or OR4 (N1795, N1790, N576, N1198, N698);
buf BUF1 (N1796, N1791);
buf BUF1 (N1797, N1769);
or OR4 (N1798, N1787, N128, N907, N177);
and AND2 (N1799, N1798, N1471);
xor XOR2 (N1800, N1781, N1719);
nand NAND2 (N1801, N1795, N930);
nor NOR4 (N1802, N1778, N1355, N593, N956);
or OR3 (N1803, N1797, N1490, N289);
buf BUF1 (N1804, N1803);
not NOT1 (N1805, N1796);
nand NAND3 (N1806, N1804, N669, N649);
nor NOR2 (N1807, N1788, N47);
nor NOR4 (N1808, N1789, N1667, N881, N845);
nor NOR2 (N1809, N1800, N485);
xor XOR2 (N1810, N1792, N117);
and AND3 (N1811, N1807, N1363, N818);
buf BUF1 (N1812, N1799);
buf BUF1 (N1813, N1805);
or OR4 (N1814, N1811, N1664, N571, N1108);
and AND3 (N1815, N1809, N872, N422);
or OR4 (N1816, N1815, N520, N1232, N80);
and AND3 (N1817, N1812, N1119, N1047);
buf BUF1 (N1818, N1814);
buf BUF1 (N1819, N1817);
buf BUF1 (N1820, N1808);
nor NOR2 (N1821, N1806, N339);
not NOT1 (N1822, N1818);
not NOT1 (N1823, N1820);
or OR3 (N1824, N1801, N92, N1803);
not NOT1 (N1825, N1813);
not NOT1 (N1826, N1810);
nand NAND2 (N1827, N1819, N487);
or OR3 (N1828, N1826, N416, N530);
or OR3 (N1829, N1816, N1580, N993);
nand NAND2 (N1830, N1822, N1062);
not NOT1 (N1831, N1828);
nor NOR2 (N1832, N1823, N1025);
xor XOR2 (N1833, N1832, N176);
buf BUF1 (N1834, N1824);
buf BUF1 (N1835, N1830);
nand NAND2 (N1836, N1821, N1636);
buf BUF1 (N1837, N1835);
and AND4 (N1838, N1794, N383, N251, N278);
xor XOR2 (N1839, N1838, N431);
and AND4 (N1840, N1825, N695, N1581, N380);
nor NOR3 (N1841, N1802, N498, N1432);
and AND2 (N1842, N1827, N93);
nand NAND2 (N1843, N1842, N1512);
or OR3 (N1844, N1829, N166, N840);
nor NOR3 (N1845, N1839, N1765, N1202);
nor NOR3 (N1846, N1841, N981, N1595);
buf BUF1 (N1847, N1831);
or OR2 (N1848, N1845, N1633);
buf BUF1 (N1849, N1847);
and AND4 (N1850, N1834, N530, N763, N765);
and AND2 (N1851, N1837, N716);
nand NAND4 (N1852, N1848, N772, N776, N1110);
xor XOR2 (N1853, N1846, N1185);
xor XOR2 (N1854, N1851, N178);
or OR3 (N1855, N1850, N1783, N231);
xor XOR2 (N1856, N1854, N1514);
not NOT1 (N1857, N1855);
nand NAND2 (N1858, N1843, N1020);
and AND4 (N1859, N1849, N1325, N707, N1212);
nor NOR2 (N1860, N1852, N310);
nand NAND4 (N1861, N1844, N1634, N901, N1144);
not NOT1 (N1862, N1836);
and AND2 (N1863, N1860, N1142);
xor XOR2 (N1864, N1863, N907);
nand NAND4 (N1865, N1862, N965, N232, N32);
buf BUF1 (N1866, N1853);
and AND2 (N1867, N1840, N538);
not NOT1 (N1868, N1861);
and AND4 (N1869, N1867, N790, N425, N413);
nand NAND2 (N1870, N1864, N26);
not NOT1 (N1871, N1857);
or OR2 (N1872, N1833, N100);
nor NOR4 (N1873, N1872, N1350, N717, N200);
nor NOR2 (N1874, N1871, N835);
or OR3 (N1875, N1865, N726, N1751);
not NOT1 (N1876, N1869);
or OR3 (N1877, N1859, N492, N61);
nand NAND4 (N1878, N1873, N768, N662, N978);
buf BUF1 (N1879, N1877);
xor XOR2 (N1880, N1866, N205);
xor XOR2 (N1881, N1879, N53);
nor NOR2 (N1882, N1876, N397);
buf BUF1 (N1883, N1874);
nand NAND2 (N1884, N1881, N552);
nand NAND3 (N1885, N1884, N1595, N1640);
not NOT1 (N1886, N1885);
nor NOR2 (N1887, N1886, N1436);
nand NAND4 (N1888, N1870, N1083, N1011, N653);
not NOT1 (N1889, N1882);
and AND2 (N1890, N1868, N726);
nor NOR4 (N1891, N1890, N1094, N862, N302);
buf BUF1 (N1892, N1880);
nand NAND2 (N1893, N1888, N1646);
xor XOR2 (N1894, N1893, N731);
nand NAND4 (N1895, N1891, N491, N835, N624);
xor XOR2 (N1896, N1858, N677);
nor NOR3 (N1897, N1875, N1042, N562);
buf BUF1 (N1898, N1856);
and AND2 (N1899, N1895, N1659);
not NOT1 (N1900, N1892);
buf BUF1 (N1901, N1894);
nor NOR3 (N1902, N1899, N1016, N1467);
nand NAND3 (N1903, N1901, N1748, N381);
xor XOR2 (N1904, N1900, N1132);
nand NAND4 (N1905, N1883, N581, N658, N1208);
and AND4 (N1906, N1897, N570, N1659, N354);
buf BUF1 (N1907, N1903);
not NOT1 (N1908, N1907);
xor XOR2 (N1909, N1889, N1899);
nor NOR4 (N1910, N1896, N476, N522, N878);
xor XOR2 (N1911, N1878, N181);
buf BUF1 (N1912, N1904);
buf BUF1 (N1913, N1911);
nor NOR4 (N1914, N1910, N1200, N1603, N1352);
and AND2 (N1915, N1912, N730);
or OR2 (N1916, N1908, N779);
nand NAND3 (N1917, N1909, N1444, N1715);
and AND2 (N1918, N1906, N635);
not NOT1 (N1919, N1898);
nand NAND3 (N1920, N1917, N401, N491);
and AND3 (N1921, N1887, N1553, N1918);
or OR4 (N1922, N764, N129, N1127, N976);
nand NAND2 (N1923, N1916, N1170);
not NOT1 (N1924, N1905);
and AND4 (N1925, N1921, N1077, N960, N1731);
nand NAND4 (N1926, N1919, N271, N1479, N1297);
nor NOR3 (N1927, N1914, N1676, N512);
or OR4 (N1928, N1927, N1888, N1857, N1914);
not NOT1 (N1929, N1913);
and AND4 (N1930, N1924, N1625, N1502, N448);
nor NOR4 (N1931, N1929, N1546, N94, N228);
buf BUF1 (N1932, N1922);
nand NAND3 (N1933, N1926, N1896, N1803);
buf BUF1 (N1934, N1933);
and AND3 (N1935, N1928, N1189, N493);
and AND3 (N1936, N1934, N531, N1572);
and AND4 (N1937, N1935, N889, N1730, N1835);
not NOT1 (N1938, N1930);
buf BUF1 (N1939, N1936);
xor XOR2 (N1940, N1925, N1062);
nor NOR2 (N1941, N1939, N964);
buf BUF1 (N1942, N1932);
not NOT1 (N1943, N1920);
not NOT1 (N1944, N1923);
buf BUF1 (N1945, N1931);
nand NAND3 (N1946, N1942, N939, N1717);
not NOT1 (N1947, N1943);
nand NAND4 (N1948, N1937, N498, N1568, N399);
nor NOR4 (N1949, N1946, N955, N1558, N1331);
buf BUF1 (N1950, N1940);
xor XOR2 (N1951, N1950, N1118);
nor NOR4 (N1952, N1902, N1123, N1153, N756);
and AND3 (N1953, N1948, N310, N1952);
or OR4 (N1954, N630, N1833, N1050, N1475);
nor NOR2 (N1955, N1949, N1844);
buf BUF1 (N1956, N1945);
xor XOR2 (N1957, N1941, N1556);
or OR4 (N1958, N1955, N751, N967, N1174);
not NOT1 (N1959, N1947);
buf BUF1 (N1960, N1958);
not NOT1 (N1961, N1938);
not NOT1 (N1962, N1953);
nand NAND2 (N1963, N1956, N473);
xor XOR2 (N1964, N1963, N712);
and AND4 (N1965, N1961, N659, N1874, N1399);
or OR3 (N1966, N1944, N207, N1166);
or OR3 (N1967, N1915, N549, N743);
not NOT1 (N1968, N1964);
or OR2 (N1969, N1959, N1425);
or OR2 (N1970, N1966, N166);
not NOT1 (N1971, N1968);
or OR3 (N1972, N1951, N1636, N326);
nand NAND4 (N1973, N1972, N873, N1326, N1958);
xor XOR2 (N1974, N1971, N1519);
not NOT1 (N1975, N1960);
not NOT1 (N1976, N1974);
nor NOR4 (N1977, N1976, N1901, N212, N1262);
xor XOR2 (N1978, N1970, N526);
xor XOR2 (N1979, N1962, N1336);
and AND2 (N1980, N1975, N1082);
buf BUF1 (N1981, N1957);
and AND4 (N1982, N1981, N1575, N1790, N816);
and AND3 (N1983, N1982, N449, N377);
nor NOR3 (N1984, N1978, N60, N1579);
nor NOR4 (N1985, N1973, N469, N1459, N1544);
and AND2 (N1986, N1969, N366);
nor NOR2 (N1987, N1983, N1162);
and AND2 (N1988, N1977, N1545);
xor XOR2 (N1989, N1980, N375);
not NOT1 (N1990, N1954);
buf BUF1 (N1991, N1967);
not NOT1 (N1992, N1965);
nand NAND3 (N1993, N1990, N1933, N1848);
not NOT1 (N1994, N1979);
nor NOR4 (N1995, N1991, N87, N1867, N1448);
not NOT1 (N1996, N1989);
nor NOR2 (N1997, N1994, N65);
or OR2 (N1998, N1988, N323);
xor XOR2 (N1999, N1984, N1398);
nand NAND2 (N2000, N1993, N866);
not NOT1 (N2001, N1999);
buf BUF1 (N2002, N1998);
buf BUF1 (N2003, N1997);
xor XOR2 (N2004, N1996, N1703);
nor NOR3 (N2005, N1992, N1946, N1939);
and AND4 (N2006, N2001, N1157, N466, N504);
nor NOR4 (N2007, N2002, N1549, N130, N268);
or OR2 (N2008, N1985, N198);
and AND2 (N2009, N1987, N885);
nor NOR3 (N2010, N2008, N1547, N233);
not NOT1 (N2011, N2010);
or OR3 (N2012, N2003, N1337, N60);
or OR2 (N2013, N2005, N1232);
nor NOR4 (N2014, N1995, N1012, N1206, N764);
or OR4 (N2015, N2004, N489, N498, N13);
nor NOR4 (N2016, N2014, N1361, N1394, N1447);
or OR4 (N2017, N2000, N141, N967, N809);
nand NAND2 (N2018, N2015, N149);
or OR2 (N2019, N2012, N268);
xor XOR2 (N2020, N1986, N97);
or OR3 (N2021, N2019, N1542, N175);
and AND4 (N2022, N2006, N11, N576, N1406);
nor NOR2 (N2023, N2009, N201);
xor XOR2 (N2024, N2011, N851);
buf BUF1 (N2025, N2007);
not NOT1 (N2026, N2018);
and AND2 (N2027, N2025, N116);
or OR4 (N2028, N2021, N650, N1121, N185);
buf BUF1 (N2029, N2026);
nand NAND3 (N2030, N2027, N1254, N18);
or OR3 (N2031, N2013, N970, N1479);
buf BUF1 (N2032, N2028);
nand NAND2 (N2033, N2032, N734);
and AND3 (N2034, N2023, N1845, N1676);
not NOT1 (N2035, N2030);
nor NOR3 (N2036, N2034, N1769, N1049);
nor NOR2 (N2037, N2029, N788);
or OR4 (N2038, N2022, N1703, N1744, N1109);
nand NAND2 (N2039, N2038, N926);
buf BUF1 (N2040, N2024);
not NOT1 (N2041, N2035);
and AND3 (N2042, N2031, N417, N1373);
and AND2 (N2043, N2016, N2004);
not NOT1 (N2044, N2043);
not NOT1 (N2045, N2042);
or OR4 (N2046, N2033, N1528, N1114, N1631);
buf BUF1 (N2047, N2020);
or OR2 (N2048, N2039, N150);
nand NAND4 (N2049, N2047, N382, N1320, N1772);
nand NAND3 (N2050, N2045, N1392, N1562);
nand NAND4 (N2051, N2041, N362, N306, N2048);
and AND4 (N2052, N625, N103, N1321, N2009);
buf BUF1 (N2053, N2049);
not NOT1 (N2054, N2036);
buf BUF1 (N2055, N2046);
buf BUF1 (N2056, N2044);
nand NAND4 (N2057, N2051, N1014, N1608, N1498);
buf BUF1 (N2058, N2052);
or OR2 (N2059, N2056, N1546);
and AND2 (N2060, N2058, N1719);
nand NAND4 (N2061, N2040, N521, N1757, N1206);
nand NAND4 (N2062, N2057, N304, N1073, N1974);
nor NOR3 (N2063, N2055, N472, N821);
nor NOR4 (N2064, N2063, N488, N1078, N998);
and AND3 (N2065, N2060, N2055, N11);
and AND3 (N2066, N2053, N220, N783);
not NOT1 (N2067, N2059);
or OR2 (N2068, N2066, N1852);
nand NAND4 (N2069, N2062, N735, N1838, N1177);
nor NOR2 (N2070, N2037, N1009);
nand NAND4 (N2071, N2061, N743, N1848, N1594);
buf BUF1 (N2072, N2054);
nand NAND4 (N2073, N2071, N146, N546, N518);
or OR3 (N2074, N2069, N809, N1365);
xor XOR2 (N2075, N2074, N2028);
buf BUF1 (N2076, N2050);
or OR4 (N2077, N2064, N509, N1864, N1346);
nand NAND3 (N2078, N2076, N260, N1066);
or OR2 (N2079, N2067, N752);
nand NAND3 (N2080, N2079, N1492, N1758);
or OR4 (N2081, N2065, N1646, N1095, N108);
nand NAND3 (N2082, N2077, N85, N1598);
not NOT1 (N2083, N2068);
and AND4 (N2084, N2070, N214, N1543, N1563);
and AND4 (N2085, N2072, N1918, N2048, N322);
and AND4 (N2086, N2078, N1023, N1181, N1334);
and AND2 (N2087, N2075, N728);
and AND4 (N2088, N2082, N1638, N174, N938);
and AND4 (N2089, N2083, N1164, N289, N1365);
and AND3 (N2090, N2085, N1462, N1314);
nand NAND3 (N2091, N2084, N105, N1569);
and AND3 (N2092, N2087, N1007, N1349);
xor XOR2 (N2093, N2017, N1778);
not NOT1 (N2094, N2073);
and AND3 (N2095, N2092, N2065, N642);
nor NOR2 (N2096, N2091, N1835);
nor NOR4 (N2097, N2096, N1625, N1638, N1556);
nor NOR3 (N2098, N2080, N809, N1190);
nand NAND3 (N2099, N2089, N551, N655);
nand NAND3 (N2100, N2094, N397, N982);
nor NOR3 (N2101, N2098, N474, N1816);
xor XOR2 (N2102, N2097, N59);
and AND2 (N2103, N2099, N1374);
xor XOR2 (N2104, N2100, N2010);
and AND3 (N2105, N2104, N558, N160);
nand NAND2 (N2106, N2095, N1320);
not NOT1 (N2107, N2103);
buf BUF1 (N2108, N2105);
and AND3 (N2109, N2090, N105, N605);
buf BUF1 (N2110, N2088);
nor NOR2 (N2111, N2086, N593);
xor XOR2 (N2112, N2107, N771);
xor XOR2 (N2113, N2081, N787);
nand NAND3 (N2114, N2106, N1671, N1264);
buf BUF1 (N2115, N2101);
buf BUF1 (N2116, N2114);
xor XOR2 (N2117, N2112, N1527);
xor XOR2 (N2118, N2109, N2102);
nor NOR4 (N2119, N1781, N1865, N289, N1934);
nand NAND2 (N2120, N2113, N433);
nand NAND4 (N2121, N2117, N400, N548, N457);
and AND3 (N2122, N2118, N84, N19);
not NOT1 (N2123, N2116);
buf BUF1 (N2124, N2108);
not NOT1 (N2125, N2124);
not NOT1 (N2126, N2123);
xor XOR2 (N2127, N2122, N1058);
and AND2 (N2128, N2093, N1565);
and AND2 (N2129, N2121, N144);
not NOT1 (N2130, N2128);
and AND4 (N2131, N2129, N1750, N1738, N150);
nand NAND3 (N2132, N2120, N1412, N1996);
not NOT1 (N2133, N2119);
buf BUF1 (N2134, N2126);
buf BUF1 (N2135, N2125);
buf BUF1 (N2136, N2131);
nor NOR2 (N2137, N2136, N1828);
nand NAND4 (N2138, N2135, N2110, N1667, N1672);
or OR3 (N2139, N114, N1970, N1152);
not NOT1 (N2140, N2132);
and AND4 (N2141, N2139, N106, N1222, N30);
or OR2 (N2142, N2137, N1314);
and AND2 (N2143, N2130, N1802);
and AND3 (N2144, N2134, N1943, N377);
not NOT1 (N2145, N2143);
nor NOR4 (N2146, N2133, N243, N930, N1427);
xor XOR2 (N2147, N2144, N2003);
nand NAND2 (N2148, N2127, N65);
xor XOR2 (N2149, N2145, N406);
and AND2 (N2150, N2147, N1540);
or OR4 (N2151, N2141, N764, N114, N784);
not NOT1 (N2152, N2149);
nand NAND3 (N2153, N2151, N959, N2051);
nand NAND2 (N2154, N2146, N574);
not NOT1 (N2155, N2140);
and AND4 (N2156, N2153, N1903, N1029, N1653);
not NOT1 (N2157, N2148);
and AND3 (N2158, N2142, N1592, N16);
xor XOR2 (N2159, N2158, N1318);
nor NOR4 (N2160, N2138, N1691, N1922, N48);
xor XOR2 (N2161, N2111, N474);
or OR4 (N2162, N2154, N1751, N870, N1151);
buf BUF1 (N2163, N2161);
and AND2 (N2164, N2155, N1738);
and AND3 (N2165, N2115, N1015, N1954);
not NOT1 (N2166, N2164);
nand NAND4 (N2167, N2156, N1321, N1634, N141);
not NOT1 (N2168, N2152);
not NOT1 (N2169, N2157);
or OR3 (N2170, N2162, N1639, N1451);
and AND3 (N2171, N2169, N1891, N1406);
xor XOR2 (N2172, N2163, N408);
or OR3 (N2173, N2165, N713, N342);
nand NAND2 (N2174, N2168, N571);
and AND3 (N2175, N2166, N352, N1501);
xor XOR2 (N2176, N2175, N297);
nand NAND4 (N2177, N2174, N35, N1029, N1003);
buf BUF1 (N2178, N2170);
nor NOR2 (N2179, N2178, N359);
nor NOR3 (N2180, N2167, N2061, N1771);
not NOT1 (N2181, N2177);
not NOT1 (N2182, N2179);
buf BUF1 (N2183, N2159);
not NOT1 (N2184, N2180);
nand NAND3 (N2185, N2181, N1649, N1562);
and AND4 (N2186, N2150, N739, N1238, N367);
nand NAND3 (N2187, N2172, N1688, N1135);
xor XOR2 (N2188, N2184, N1331);
or OR3 (N2189, N2186, N681, N1556);
nor NOR4 (N2190, N2187, N1950, N1740, N458);
or OR2 (N2191, N2171, N730);
and AND4 (N2192, N2190, N331, N1078, N1194);
nand NAND3 (N2193, N2192, N1727, N837);
nor NOR2 (N2194, N2191, N2090);
nand NAND2 (N2195, N2183, N132);
not NOT1 (N2196, N2182);
not NOT1 (N2197, N2195);
or OR2 (N2198, N2194, N822);
nand NAND2 (N2199, N2189, N291);
buf BUF1 (N2200, N2193);
xor XOR2 (N2201, N2199, N1309);
buf BUF1 (N2202, N2160);
nand NAND3 (N2203, N2198, N300, N993);
xor XOR2 (N2204, N2203, N638);
xor XOR2 (N2205, N2185, N1468);
nor NOR3 (N2206, N2200, N627, N391);
nand NAND4 (N2207, N2204, N780, N1244, N964);
nand NAND2 (N2208, N2202, N964);
xor XOR2 (N2209, N2196, N1821);
not NOT1 (N2210, N2201);
nand NAND4 (N2211, N2173, N171, N1007, N1481);
not NOT1 (N2212, N2197);
xor XOR2 (N2213, N2209, N1829);
not NOT1 (N2214, N2205);
not NOT1 (N2215, N2188);
buf BUF1 (N2216, N2211);
xor XOR2 (N2217, N2208, N1912);
buf BUF1 (N2218, N2216);
nor NOR2 (N2219, N2214, N797);
buf BUF1 (N2220, N2217);
and AND3 (N2221, N2215, N117, N362);
and AND2 (N2222, N2212, N684);
nand NAND4 (N2223, N2220, N2078, N234, N1092);
not NOT1 (N2224, N2223);
buf BUF1 (N2225, N2222);
and AND2 (N2226, N2210, N1606);
nor NOR3 (N2227, N2207, N698, N1890);
or OR3 (N2228, N2225, N1166, N2169);
nor NOR3 (N2229, N2221, N739, N375);
buf BUF1 (N2230, N2219);
nand NAND3 (N2231, N2227, N1294, N2131);
and AND2 (N2232, N2231, N270);
not NOT1 (N2233, N2229);
nand NAND3 (N2234, N2176, N1603, N1644);
nand NAND2 (N2235, N2224, N315);
and AND2 (N2236, N2228, N439);
buf BUF1 (N2237, N2233);
or OR2 (N2238, N2230, N1739);
nand NAND3 (N2239, N2232, N1674, N837);
or OR4 (N2240, N2206, N831, N59, N817);
not NOT1 (N2241, N2226);
buf BUF1 (N2242, N2234);
or OR2 (N2243, N2235, N1447);
buf BUF1 (N2244, N2242);
nor NOR4 (N2245, N2243, N706, N2243, N1440);
and AND2 (N2246, N2241, N888);
xor XOR2 (N2247, N2236, N471);
nand NAND4 (N2248, N2239, N108, N30, N935);
xor XOR2 (N2249, N2238, N2038);
xor XOR2 (N2250, N2240, N1018);
not NOT1 (N2251, N2213);
not NOT1 (N2252, N2248);
or OR4 (N2253, N2247, N1837, N1835, N2114);
nor NOR3 (N2254, N2237, N1770, N362);
not NOT1 (N2255, N2249);
nor NOR2 (N2256, N2250, N873);
not NOT1 (N2257, N2254);
or OR4 (N2258, N2251, N2121, N1675, N957);
or OR2 (N2259, N2218, N1091);
and AND3 (N2260, N2246, N1470, N745);
nor NOR3 (N2261, N2258, N1692, N2145);
or OR2 (N2262, N2260, N1921);
and AND2 (N2263, N2244, N117);
nand NAND3 (N2264, N2255, N174, N1281);
not NOT1 (N2265, N2245);
not NOT1 (N2266, N2264);
and AND3 (N2267, N2253, N1728, N500);
and AND3 (N2268, N2265, N2180, N1785);
not NOT1 (N2269, N2261);
nor NOR4 (N2270, N2262, N1254, N1838, N2222);
nand NAND2 (N2271, N2257, N2065);
not NOT1 (N2272, N2269);
or OR3 (N2273, N2266, N1855, N61);
nor NOR2 (N2274, N2263, N1506);
or OR2 (N2275, N2259, N984);
and AND4 (N2276, N2267, N510, N2256, N747);
and AND3 (N2277, N1490, N745, N1705);
not NOT1 (N2278, N2271);
buf BUF1 (N2279, N2272);
buf BUF1 (N2280, N2268);
or OR4 (N2281, N2275, N1772, N1356, N1603);
and AND4 (N2282, N2252, N1135, N2220, N2161);
or OR4 (N2283, N2274, N1693, N1729, N1680);
or OR3 (N2284, N2283, N394, N566);
and AND2 (N2285, N2280, N152);
and AND2 (N2286, N2281, N332);
nor NOR3 (N2287, N2276, N1869, N182);
or OR4 (N2288, N2284, N263, N297, N2074);
nor NOR2 (N2289, N2278, N1089);
or OR3 (N2290, N2286, N273, N1020);
xor XOR2 (N2291, N2290, N2287);
not NOT1 (N2292, N509);
nand NAND3 (N2293, N2292, N732, N519);
not NOT1 (N2294, N2273);
or OR4 (N2295, N2282, N1974, N652, N176);
buf BUF1 (N2296, N2289);
or OR3 (N2297, N2277, N727, N1491);
nand NAND2 (N2298, N2285, N1377);
xor XOR2 (N2299, N2291, N1869);
or OR2 (N2300, N2297, N1099);
or OR3 (N2301, N2279, N1062, N1284);
xor XOR2 (N2302, N2299, N1091);
nand NAND4 (N2303, N2296, N1620, N1864, N2153);
or OR4 (N2304, N2302, N2056, N259, N2195);
xor XOR2 (N2305, N2298, N876);
nand NAND4 (N2306, N2304, N2264, N745, N1307);
not NOT1 (N2307, N2300);
nor NOR3 (N2308, N2288, N599, N2000);
not NOT1 (N2309, N2295);
xor XOR2 (N2310, N2309, N933);
nor NOR4 (N2311, N2301, N870, N867, N1030);
xor XOR2 (N2312, N2308, N203);
xor XOR2 (N2313, N2306, N175);
not NOT1 (N2314, N2293);
or OR2 (N2315, N2294, N120);
nand NAND2 (N2316, N2307, N1101);
nand NAND2 (N2317, N2312, N375);
or OR3 (N2318, N2316, N776, N240);
nand NAND3 (N2319, N2314, N1166, N413);
buf BUF1 (N2320, N2319);
buf BUF1 (N2321, N2305);
xor XOR2 (N2322, N2311, N1847);
or OR3 (N2323, N2310, N1449, N2221);
xor XOR2 (N2324, N2322, N332);
nor NOR3 (N2325, N2270, N466, N565);
nor NOR4 (N2326, N2320, N2273, N1037, N854);
xor XOR2 (N2327, N2326, N1513);
buf BUF1 (N2328, N2313);
nand NAND4 (N2329, N2325, N1224, N4, N1940);
and AND3 (N2330, N2315, N1031, N2301);
and AND2 (N2331, N2330, N2035);
or OR3 (N2332, N2328, N2269, N1369);
not NOT1 (N2333, N2331);
nand NAND2 (N2334, N2327, N1293);
buf BUF1 (N2335, N2324);
nand NAND2 (N2336, N2333, N1896);
and AND4 (N2337, N2332, N231, N2213, N1569);
nand NAND2 (N2338, N2337, N793);
xor XOR2 (N2339, N2323, N1610);
nor NOR4 (N2340, N2334, N1035, N1522, N1773);
and AND4 (N2341, N2303, N332, N935, N807);
xor XOR2 (N2342, N2341, N1163);
nor NOR3 (N2343, N2317, N1185, N1845);
buf BUF1 (N2344, N2342);
and AND3 (N2345, N2335, N1177, N1364);
nand NAND3 (N2346, N2340, N83, N163);
or OR3 (N2347, N2339, N979, N1242);
xor XOR2 (N2348, N2329, N845);
buf BUF1 (N2349, N2343);
not NOT1 (N2350, N2347);
buf BUF1 (N2351, N2346);
nor NOR2 (N2352, N2344, N90);
not NOT1 (N2353, N2352);
not NOT1 (N2354, N2349);
not NOT1 (N2355, N2351);
xor XOR2 (N2356, N2353, N1885);
xor XOR2 (N2357, N2355, N1248);
buf BUF1 (N2358, N2345);
nand NAND3 (N2359, N2354, N1986, N207);
not NOT1 (N2360, N2348);
nor NOR3 (N2361, N2321, N799, N1694);
nand NAND4 (N2362, N2338, N1448, N1435, N1921);
not NOT1 (N2363, N2360);
nand NAND2 (N2364, N2357, N1439);
nor NOR2 (N2365, N2318, N493);
buf BUF1 (N2366, N2336);
nor NOR4 (N2367, N2366, N1737, N1203, N1421);
not NOT1 (N2368, N2350);
nor NOR3 (N2369, N2363, N463, N1382);
buf BUF1 (N2370, N2365);
nor NOR3 (N2371, N2368, N2204, N2085);
nor NOR4 (N2372, N2358, N668, N337, N556);
nand NAND2 (N2373, N2361, N389);
and AND4 (N2374, N2370, N287, N1419, N568);
nor NOR4 (N2375, N2372, N523, N2100, N2178);
nor NOR3 (N2376, N2375, N293, N1550);
xor XOR2 (N2377, N2371, N1453);
and AND4 (N2378, N2373, N725, N590, N1529);
xor XOR2 (N2379, N2364, N1320);
buf BUF1 (N2380, N2369);
or OR2 (N2381, N2374, N681);
xor XOR2 (N2382, N2381, N1272);
not NOT1 (N2383, N2359);
or OR3 (N2384, N2380, N498, N1489);
or OR4 (N2385, N2379, N1707, N1411, N1322);
xor XOR2 (N2386, N2382, N640);
buf BUF1 (N2387, N2376);
and AND2 (N2388, N2362, N1098);
and AND4 (N2389, N2385, N2142, N517, N2218);
and AND3 (N2390, N2389, N1160, N884);
nand NAND3 (N2391, N2356, N2058, N15);
nand NAND4 (N2392, N2387, N1256, N741, N1020);
xor XOR2 (N2393, N2378, N844);
not NOT1 (N2394, N2392);
xor XOR2 (N2395, N2390, N1745);
nor NOR4 (N2396, N2386, N663, N477, N1555);
or OR4 (N2397, N2367, N2209, N321, N1521);
nor NOR2 (N2398, N2393, N562);
not NOT1 (N2399, N2377);
and AND3 (N2400, N2396, N1478, N1408);
buf BUF1 (N2401, N2383);
nor NOR3 (N2402, N2388, N1671, N1970);
not NOT1 (N2403, N2400);
buf BUF1 (N2404, N2394);
nor NOR2 (N2405, N2391, N887);
and AND3 (N2406, N2397, N1677, N1717);
xor XOR2 (N2407, N2405, N1925);
xor XOR2 (N2408, N2398, N2360);
or OR2 (N2409, N2403, N2373);
nand NAND3 (N2410, N2384, N1899, N1637);
and AND3 (N2411, N2406, N406, N1858);
buf BUF1 (N2412, N2399);
xor XOR2 (N2413, N2409, N1503);
not NOT1 (N2414, N2402);
not NOT1 (N2415, N2408);
nor NOR2 (N2416, N2411, N1730);
nand NAND4 (N2417, N2395, N2282, N54, N2335);
not NOT1 (N2418, N2401);
not NOT1 (N2419, N2414);
nor NOR4 (N2420, N2412, N1044, N2010, N1015);
and AND4 (N2421, N2418, N149, N749, N2379);
buf BUF1 (N2422, N2410);
nand NAND2 (N2423, N2413, N2404);
not NOT1 (N2424, N1040);
nor NOR2 (N2425, N2422, N2017);
nor NOR4 (N2426, N2421, N1820, N1988, N2401);
nor NOR4 (N2427, N2407, N1285, N92, N222);
buf BUF1 (N2428, N2416);
and AND3 (N2429, N2427, N1529, N2351);
nor NOR2 (N2430, N2425, N2052);
nand NAND2 (N2431, N2419, N839);
not NOT1 (N2432, N2424);
nor NOR2 (N2433, N2431, N1736);
xor XOR2 (N2434, N2433, N459);
nand NAND3 (N2435, N2417, N585, N2110);
nand NAND2 (N2436, N2415, N2317);
and AND4 (N2437, N2426, N1596, N1013, N2208);
and AND4 (N2438, N2428, N434, N1271, N759);
or OR3 (N2439, N2432, N1074, N765);
not NOT1 (N2440, N2437);
or OR2 (N2441, N2440, N741);
and AND2 (N2442, N2439, N610);
or OR4 (N2443, N2420, N2215, N1443, N1809);
nand NAND2 (N2444, N2435, N2246);
nand NAND4 (N2445, N2430, N2109, N2040, N2183);
nor NOR2 (N2446, N2429, N1952);
and AND2 (N2447, N2445, N555);
xor XOR2 (N2448, N2436, N1001);
buf BUF1 (N2449, N2441);
xor XOR2 (N2450, N2434, N569);
and AND2 (N2451, N2449, N656);
nor NOR4 (N2452, N2443, N177, N2048, N1889);
or OR4 (N2453, N2438, N2412, N1686, N395);
xor XOR2 (N2454, N2453, N2377);
buf BUF1 (N2455, N2450);
nor NOR3 (N2456, N2451, N1118, N2013);
not NOT1 (N2457, N2423);
buf BUF1 (N2458, N2444);
nor NOR2 (N2459, N2448, N141);
nand NAND2 (N2460, N2446, N812);
nand NAND4 (N2461, N2442, N1669, N241, N1695);
nand NAND3 (N2462, N2452, N1406, N1812);
nor NOR2 (N2463, N2462, N1073);
nor NOR3 (N2464, N2458, N1764, N339);
nand NAND3 (N2465, N2460, N266, N2371);
nor NOR2 (N2466, N2454, N535);
and AND4 (N2467, N2447, N1186, N2201, N1515);
xor XOR2 (N2468, N2456, N143);
or OR3 (N2469, N2463, N1145, N99);
xor XOR2 (N2470, N2464, N394);
nor NOR4 (N2471, N2465, N1561, N2123, N1767);
not NOT1 (N2472, N2470);
xor XOR2 (N2473, N2467, N450);
buf BUF1 (N2474, N2459);
buf BUF1 (N2475, N2466);
buf BUF1 (N2476, N2471);
nor NOR3 (N2477, N2475, N9, N238);
xor XOR2 (N2478, N2461, N592);
nand NAND2 (N2479, N2455, N2);
nor NOR4 (N2480, N2473, N1665, N153, N1694);
nor NOR2 (N2481, N2476, N1204);
or OR3 (N2482, N2479, N161, N1069);
and AND3 (N2483, N2477, N27, N2378);
xor XOR2 (N2484, N2482, N1843);
and AND3 (N2485, N2484, N2092, N1640);
nand NAND3 (N2486, N2474, N1002, N196);
xor XOR2 (N2487, N2468, N1665);
nand NAND4 (N2488, N2483, N2244, N2069, N1602);
nor NOR2 (N2489, N2480, N2385);
nor NOR4 (N2490, N2472, N2037, N117, N2084);
or OR2 (N2491, N2487, N233);
and AND2 (N2492, N2491, N1356);
nand NAND3 (N2493, N2469, N1267, N467);
nor NOR3 (N2494, N2493, N1061, N773);
not NOT1 (N2495, N2494);
not NOT1 (N2496, N2492);
and AND2 (N2497, N2488, N1431);
nand NAND3 (N2498, N2497, N256, N2143);
and AND3 (N2499, N2495, N1712, N2055);
nand NAND2 (N2500, N2485, N715);
buf BUF1 (N2501, N2457);
or OR4 (N2502, N2490, N1900, N1238, N1022);
xor XOR2 (N2503, N2489, N668);
nor NOR3 (N2504, N2501, N1898, N964);
not NOT1 (N2505, N2502);
xor XOR2 (N2506, N2504, N336);
not NOT1 (N2507, N2506);
nor NOR3 (N2508, N2486, N80, N856);
nor NOR3 (N2509, N2507, N105, N321);
nor NOR2 (N2510, N2509, N334);
buf BUF1 (N2511, N2498);
or OR2 (N2512, N2505, N801);
xor XOR2 (N2513, N2511, N2181);
endmodule