// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19;

output N506,N516,N510,N517,N518,N514,N515,N512,N498,N519;

not NOT1 (N20, N2);
xor XOR2 (N21, N5, N4);
not NOT1 (N22, N19);
not NOT1 (N23, N18);
or OR3 (N24, N16, N23, N15);
nor NOR4 (N25, N6, N3, N16, N9);
buf BUF1 (N26, N23);
and AND4 (N27, N11, N10, N8, N26);
and AND4 (N28, N26, N23, N13, N23);
buf BUF1 (N29, N6);
or OR4 (N30, N25, N5, N13, N21);
nor NOR2 (N31, N26, N1);
or OR2 (N32, N24, N10);
not NOT1 (N33, N22);
not NOT1 (N34, N14);
and AND3 (N35, N26, N2, N28);
buf BUF1 (N36, N29);
xor XOR2 (N37, N22, N8);
buf BUF1 (N38, N20);
xor XOR2 (N39, N34, N18);
or OR2 (N40, N37, N11);
xor XOR2 (N41, N30, N34);
xor XOR2 (N42, N35, N33);
and AND4 (N43, N7, N35, N24, N26);
nor NOR3 (N44, N27, N9, N19);
buf BUF1 (N45, N32);
or OR2 (N46, N42, N38);
and AND4 (N47, N43, N38, N17, N32);
and AND4 (N48, N44, N19, N36, N38);
or OR4 (N49, N19, N31, N34, N10);
and AND2 (N50, N16, N49);
not NOT1 (N51, N32);
nor NOR4 (N52, N4, N1, N49, N17);
not NOT1 (N53, N41);
not NOT1 (N54, N47);
xor XOR2 (N55, N46, N13);
or OR2 (N56, N54, N51);
buf BUF1 (N57, N48);
buf BUF1 (N58, N31);
and AND3 (N59, N39, N39, N17);
or OR4 (N60, N56, N25, N40, N49);
or OR2 (N61, N56, N18);
and AND3 (N62, N53, N26, N4);
not NOT1 (N63, N55);
and AND4 (N64, N50, N19, N13, N40);
nor NOR2 (N65, N62, N54);
xor XOR2 (N66, N52, N15);
nand NAND2 (N67, N61, N16);
or OR3 (N68, N60, N32, N14);
xor XOR2 (N69, N66, N14);
and AND2 (N70, N58, N42);
and AND2 (N71, N64, N14);
xor XOR2 (N72, N67, N49);
nand NAND3 (N73, N70, N67, N40);
xor XOR2 (N74, N71, N53);
and AND2 (N75, N69, N46);
buf BUF1 (N76, N68);
xor XOR2 (N77, N72, N33);
not NOT1 (N78, N75);
or OR4 (N79, N74, N31, N33, N27);
not NOT1 (N80, N59);
not NOT1 (N81, N80);
or OR3 (N82, N45, N1, N16);
xor XOR2 (N83, N73, N15);
or OR3 (N84, N77, N48, N39);
not NOT1 (N85, N65);
xor XOR2 (N86, N85, N18);
or OR3 (N87, N63, N80, N52);
not NOT1 (N88, N87);
nor NOR4 (N89, N79, N63, N74, N31);
buf BUF1 (N90, N84);
buf BUF1 (N91, N82);
or OR2 (N92, N89, N19);
xor XOR2 (N93, N76, N87);
xor XOR2 (N94, N86, N10);
and AND2 (N95, N94, N37);
not NOT1 (N96, N95);
xor XOR2 (N97, N88, N75);
buf BUF1 (N98, N78);
or OR2 (N99, N81, N71);
buf BUF1 (N100, N98);
not NOT1 (N101, N100);
nor NOR4 (N102, N90, N56, N65, N63);
nand NAND2 (N103, N57, N78);
or OR4 (N104, N91, N84, N66, N23);
xor XOR2 (N105, N99, N48);
nand NAND2 (N106, N104, N46);
buf BUF1 (N107, N106);
nand NAND3 (N108, N107, N105, N77);
nor NOR4 (N109, N103, N75, N26, N16);
and AND4 (N110, N8, N12, N96, N4);
or OR4 (N111, N58, N52, N80, N69);
buf BUF1 (N112, N97);
xor XOR2 (N113, N109, N37);
xor XOR2 (N114, N110, N110);
and AND3 (N115, N113, N8, N46);
buf BUF1 (N116, N92);
not NOT1 (N117, N101);
and AND3 (N118, N108, N70, N26);
nand NAND4 (N119, N116, N13, N97, N42);
and AND4 (N120, N83, N84, N103, N102);
and AND4 (N121, N70, N61, N3, N20);
nand NAND3 (N122, N121, N76, N88);
xor XOR2 (N123, N119, N33);
buf BUF1 (N124, N93);
xor XOR2 (N125, N122, N122);
nand NAND2 (N126, N115, N56);
nor NOR4 (N127, N114, N46, N117, N85);
and AND2 (N128, N95, N69);
and AND3 (N129, N125, N10, N28);
nand NAND4 (N130, N126, N51, N38, N110);
buf BUF1 (N131, N130);
or OR4 (N132, N118, N121, N61, N71);
nand NAND2 (N133, N124, N123);
not NOT1 (N134, N126);
nor NOR2 (N135, N131, N6);
xor XOR2 (N136, N134, N94);
not NOT1 (N137, N111);
nor NOR4 (N138, N112, N36, N126, N11);
xor XOR2 (N139, N127, N93);
buf BUF1 (N140, N132);
and AND4 (N141, N137, N32, N135, N52);
nor NOR2 (N142, N10, N25);
and AND4 (N143, N136, N107, N61, N51);
or OR2 (N144, N128, N16);
not NOT1 (N145, N140);
xor XOR2 (N146, N144, N97);
and AND2 (N147, N145, N7);
or OR4 (N148, N129, N43, N92, N106);
nand NAND3 (N149, N120, N97, N17);
or OR2 (N150, N139, N45);
and AND2 (N151, N142, N102);
not NOT1 (N152, N146);
nand NAND3 (N153, N143, N8, N145);
buf BUF1 (N154, N152);
nand NAND3 (N155, N154, N132, N97);
buf BUF1 (N156, N148);
xor XOR2 (N157, N138, N120);
nor NOR2 (N158, N147, N59);
nand NAND3 (N159, N133, N117, N61);
nand NAND4 (N160, N153, N154, N148, N85);
xor XOR2 (N161, N158, N71);
not NOT1 (N162, N159);
or OR2 (N163, N151, N106);
nand NAND2 (N164, N149, N92);
nor NOR4 (N165, N161, N141, N110, N148);
nand NAND3 (N166, N127, N17, N84);
nand NAND4 (N167, N160, N142, N108, N74);
or OR4 (N168, N150, N167, N9, N88);
not NOT1 (N169, N3);
nand NAND3 (N170, N162, N71, N135);
nand NAND3 (N171, N164, N115, N102);
nor NOR4 (N172, N169, N37, N96, N126);
buf BUF1 (N173, N166);
xor XOR2 (N174, N165, N44);
xor XOR2 (N175, N155, N31);
nand NAND3 (N176, N175, N127, N91);
nor NOR3 (N177, N174, N94, N159);
nand NAND3 (N178, N168, N43, N47);
and AND3 (N179, N171, N46, N17);
buf BUF1 (N180, N173);
or OR2 (N181, N170, N122);
xor XOR2 (N182, N180, N142);
or OR3 (N183, N156, N33, N15);
nor NOR4 (N184, N172, N21, N35, N124);
nand NAND2 (N185, N181, N6);
nand NAND4 (N186, N163, N111, N23, N152);
and AND3 (N187, N185, N10, N111);
nand NAND3 (N188, N179, N144, N100);
nor NOR3 (N189, N178, N30, N148);
or OR4 (N190, N177, N84, N142, N147);
xor XOR2 (N191, N189, N59);
and AND4 (N192, N186, N108, N175, N42);
nor NOR3 (N193, N188, N178, N142);
nand NAND3 (N194, N192, N56, N156);
buf BUF1 (N195, N194);
or OR4 (N196, N157, N126, N34, N121);
buf BUF1 (N197, N183);
nand NAND2 (N198, N187, N82);
and AND4 (N199, N193, N84, N197, N171);
xor XOR2 (N200, N142, N93);
nand NAND4 (N201, N182, N184, N85, N114);
buf BUF1 (N202, N139);
not NOT1 (N203, N201);
or OR4 (N204, N196, N46, N96, N26);
nor NOR2 (N205, N202, N189);
and AND4 (N206, N191, N148, N183, N197);
nor NOR3 (N207, N204, N40, N28);
nor NOR4 (N208, N195, N100, N192, N23);
buf BUF1 (N209, N203);
nor NOR3 (N210, N205, N192, N36);
and AND3 (N211, N208, N78, N195);
nand NAND2 (N212, N190, N77);
nand NAND3 (N213, N176, N197, N25);
xor XOR2 (N214, N211, N12);
buf BUF1 (N215, N199);
buf BUF1 (N216, N209);
and AND2 (N217, N213, N39);
buf BUF1 (N218, N200);
nor NOR2 (N219, N215, N52);
or OR3 (N220, N210, N183, N129);
nor NOR3 (N221, N198, N87, N92);
and AND3 (N222, N220, N96, N30);
xor XOR2 (N223, N218, N124);
nor NOR4 (N224, N207, N135, N166, N202);
nor NOR2 (N225, N223, N80);
buf BUF1 (N226, N224);
nand NAND3 (N227, N225, N118, N129);
xor XOR2 (N228, N216, N157);
buf BUF1 (N229, N212);
nand NAND2 (N230, N219, N93);
xor XOR2 (N231, N206, N195);
buf BUF1 (N232, N214);
and AND4 (N233, N228, N72, N230, N153);
and AND3 (N234, N151, N196, N202);
nor NOR4 (N235, N231, N180, N233, N5);
nor NOR2 (N236, N102, N70);
xor XOR2 (N237, N221, N186);
or OR2 (N238, N222, N220);
buf BUF1 (N239, N237);
xor XOR2 (N240, N226, N196);
buf BUF1 (N241, N232);
nor NOR4 (N242, N229, N191, N141, N37);
not NOT1 (N243, N235);
xor XOR2 (N244, N240, N197);
not NOT1 (N245, N242);
and AND4 (N246, N239, N85, N172, N187);
nor NOR4 (N247, N245, N226, N86, N225);
not NOT1 (N248, N236);
not NOT1 (N249, N246);
nor NOR4 (N250, N248, N143, N242, N135);
and AND3 (N251, N217, N100, N147);
xor XOR2 (N252, N250, N96);
and AND4 (N253, N247, N43, N166, N3);
nor NOR2 (N254, N249, N243);
xor XOR2 (N255, N179, N18);
nand NAND3 (N256, N255, N216, N168);
buf BUF1 (N257, N256);
or OR4 (N258, N234, N93, N78, N36);
or OR4 (N259, N257, N212, N89, N190);
nand NAND2 (N260, N227, N27);
or OR3 (N261, N258, N259, N114);
xor XOR2 (N262, N192, N233);
nand NAND2 (N263, N262, N43);
nand NAND2 (N264, N254, N27);
xor XOR2 (N265, N263, N58);
not NOT1 (N266, N253);
nor NOR2 (N267, N252, N6);
not NOT1 (N268, N264);
xor XOR2 (N269, N241, N149);
nand NAND2 (N270, N251, N135);
or OR4 (N271, N266, N246, N191, N145);
and AND2 (N272, N238, N250);
buf BUF1 (N273, N269);
nand NAND4 (N274, N261, N5, N26, N256);
nand NAND3 (N275, N265, N63, N273);
not NOT1 (N276, N170);
not NOT1 (N277, N275);
and AND2 (N278, N268, N97);
and AND2 (N279, N272, N77);
buf BUF1 (N280, N270);
xor XOR2 (N281, N277, N5);
nor NOR2 (N282, N267, N140);
and AND3 (N283, N274, N149, N142);
or OR3 (N284, N281, N180, N97);
xor XOR2 (N285, N260, N83);
and AND2 (N286, N280, N205);
buf BUF1 (N287, N271);
and AND3 (N288, N287, N42, N96);
nand NAND4 (N289, N278, N218, N145, N130);
and AND2 (N290, N276, N249);
nand NAND3 (N291, N289, N54, N104);
and AND4 (N292, N286, N43, N107, N18);
or OR2 (N293, N284, N248);
not NOT1 (N294, N282);
nand NAND3 (N295, N290, N191, N4);
buf BUF1 (N296, N244);
and AND3 (N297, N283, N79, N10);
or OR2 (N298, N295, N254);
or OR2 (N299, N296, N99);
and AND3 (N300, N299, N281, N245);
not NOT1 (N301, N297);
not NOT1 (N302, N279);
buf BUF1 (N303, N301);
xor XOR2 (N304, N288, N89);
nand NAND3 (N305, N285, N165, N1);
xor XOR2 (N306, N291, N242);
and AND3 (N307, N300, N229, N49);
buf BUF1 (N308, N303);
and AND2 (N309, N308, N123);
not NOT1 (N310, N302);
nand NAND4 (N311, N304, N224, N59, N54);
and AND3 (N312, N309, N80, N162);
and AND4 (N313, N298, N69, N184, N275);
buf BUF1 (N314, N292);
nand NAND2 (N315, N311, N106);
not NOT1 (N316, N310);
buf BUF1 (N317, N312);
and AND2 (N318, N317, N227);
nor NOR4 (N319, N306, N242, N238, N94);
and AND3 (N320, N307, N24, N226);
nor NOR3 (N321, N313, N230, N221);
and AND4 (N322, N314, N120, N307, N79);
and AND4 (N323, N316, N211, N101, N91);
xor XOR2 (N324, N318, N128);
nor NOR4 (N325, N319, N254, N311, N298);
nand NAND2 (N326, N321, N58);
not NOT1 (N327, N324);
buf BUF1 (N328, N315);
nand NAND2 (N329, N322, N79);
nand NAND2 (N330, N325, N279);
or OR2 (N331, N293, N181);
buf BUF1 (N332, N305);
nor NOR4 (N333, N331, N204, N113, N313);
or OR4 (N334, N323, N329, N249, N216);
nand NAND4 (N335, N7, N70, N1, N59);
nor NOR3 (N336, N328, N105, N260);
xor XOR2 (N337, N336, N237);
buf BUF1 (N338, N330);
and AND3 (N339, N326, N112, N233);
buf BUF1 (N340, N327);
nor NOR2 (N341, N338, N234);
nor NOR2 (N342, N339, N146);
nor NOR2 (N343, N294, N95);
nand NAND3 (N344, N343, N288, N301);
or OR2 (N345, N332, N32);
nor NOR3 (N346, N334, N55, N198);
xor XOR2 (N347, N342, N340);
nor NOR4 (N348, N203, N17, N143, N278);
nor NOR4 (N349, N347, N323, N212, N274);
not NOT1 (N350, N346);
nor NOR3 (N351, N344, N286, N152);
nor NOR4 (N352, N345, N249, N283, N249);
xor XOR2 (N353, N348, N112);
xor XOR2 (N354, N349, N333);
buf BUF1 (N355, N159);
or OR3 (N356, N352, N31, N14);
not NOT1 (N357, N350);
not NOT1 (N358, N320);
not NOT1 (N359, N356);
not NOT1 (N360, N337);
not NOT1 (N361, N358);
nor NOR2 (N362, N355, N207);
and AND4 (N363, N361, N136, N279, N142);
not NOT1 (N364, N359);
xor XOR2 (N365, N363, N69);
and AND4 (N366, N360, N190, N36, N110);
not NOT1 (N367, N362);
or OR3 (N368, N365, N102, N242);
or OR4 (N369, N364, N280, N111, N327);
not NOT1 (N370, N366);
not NOT1 (N371, N354);
not NOT1 (N372, N367);
xor XOR2 (N373, N371, N210);
nand NAND3 (N374, N369, N302, N145);
and AND4 (N375, N351, N34, N295, N162);
nor NOR3 (N376, N335, N86, N196);
nor NOR4 (N377, N375, N233, N100, N221);
buf BUF1 (N378, N373);
xor XOR2 (N379, N368, N59);
and AND3 (N380, N357, N353, N189);
and AND2 (N381, N262, N269);
not NOT1 (N382, N376);
nand NAND2 (N383, N382, N354);
nor NOR2 (N384, N379, N139);
buf BUF1 (N385, N380);
and AND2 (N386, N377, N266);
buf BUF1 (N387, N383);
nor NOR2 (N388, N381, N103);
and AND4 (N389, N387, N158, N370, N26);
not NOT1 (N390, N357);
buf BUF1 (N391, N372);
xor XOR2 (N392, N385, N46);
not NOT1 (N393, N386);
or OR2 (N394, N391, N132);
and AND2 (N395, N388, N165);
nor NOR4 (N396, N384, N126, N172, N116);
or OR2 (N397, N378, N170);
nor NOR3 (N398, N341, N94, N301);
nand NAND2 (N399, N395, N82);
nand NAND2 (N400, N392, N325);
xor XOR2 (N401, N374, N63);
xor XOR2 (N402, N390, N389);
xor XOR2 (N403, N153, N19);
and AND4 (N404, N393, N174, N400, N343);
and AND2 (N405, N7, N303);
nand NAND2 (N406, N398, N59);
not NOT1 (N407, N394);
xor XOR2 (N408, N397, N50);
xor XOR2 (N409, N407, N79);
or OR4 (N410, N406, N380, N80, N362);
nor NOR2 (N411, N403, N370);
buf BUF1 (N412, N405);
nand NAND2 (N413, N408, N212);
and AND3 (N414, N411, N68, N372);
and AND2 (N415, N399, N7);
nor NOR3 (N416, N409, N17, N243);
not NOT1 (N417, N401);
or OR2 (N418, N413, N116);
nor NOR4 (N419, N402, N106, N406, N261);
buf BUF1 (N420, N414);
buf BUF1 (N421, N418);
nor NOR4 (N422, N420, N417, N325, N410);
nand NAND3 (N423, N70, N142, N270);
xor XOR2 (N424, N16, N44);
xor XOR2 (N425, N421, N277);
nand NAND2 (N426, N415, N128);
and AND2 (N427, N424, N34);
xor XOR2 (N428, N404, N123);
xor XOR2 (N429, N412, N82);
nand NAND3 (N430, N426, N188, N43);
or OR3 (N431, N429, N146, N258);
xor XOR2 (N432, N427, N107);
not NOT1 (N433, N416);
and AND2 (N434, N432, N1);
buf BUF1 (N435, N433);
nor NOR2 (N436, N425, N17);
xor XOR2 (N437, N428, N371);
or OR4 (N438, N431, N78, N196, N245);
not NOT1 (N439, N430);
buf BUF1 (N440, N419);
not NOT1 (N441, N439);
nand NAND3 (N442, N440, N63, N68);
nand NAND3 (N443, N435, N223, N231);
buf BUF1 (N444, N434);
not NOT1 (N445, N396);
or OR4 (N446, N445, N397, N121, N151);
xor XOR2 (N447, N446, N211);
nand NAND4 (N448, N422, N66, N95, N396);
and AND2 (N449, N442, N188);
and AND3 (N450, N423, N134, N156);
buf BUF1 (N451, N437);
xor XOR2 (N452, N441, N46);
or OR2 (N453, N447, N221);
nor NOR2 (N454, N451, N106);
xor XOR2 (N455, N444, N421);
not NOT1 (N456, N448);
buf BUF1 (N457, N438);
or OR4 (N458, N453, N437, N233, N339);
or OR3 (N459, N457, N242, N442);
nor NOR2 (N460, N456, N28);
nand NAND2 (N461, N443, N5);
buf BUF1 (N462, N450);
or OR4 (N463, N455, N136, N420, N152);
buf BUF1 (N464, N459);
or OR3 (N465, N461, N179, N75);
buf BUF1 (N466, N458);
nor NOR3 (N467, N452, N412, N188);
not NOT1 (N468, N460);
xor XOR2 (N469, N463, N185);
and AND4 (N470, N466, N398, N230, N162);
buf BUF1 (N471, N454);
xor XOR2 (N472, N471, N375);
or OR4 (N473, N449, N408, N266, N384);
and AND4 (N474, N467, N89, N370, N108);
buf BUF1 (N475, N462);
or OR3 (N476, N469, N32, N66);
nor NOR3 (N477, N468, N343, N400);
not NOT1 (N478, N464);
buf BUF1 (N479, N470);
and AND4 (N480, N478, N397, N388, N152);
nand NAND3 (N481, N473, N466, N236);
nor NOR4 (N482, N465, N459, N121, N331);
nand NAND2 (N483, N479, N407);
and AND3 (N484, N476, N247, N192);
not NOT1 (N485, N481);
buf BUF1 (N486, N436);
nor NOR2 (N487, N472, N164);
not NOT1 (N488, N474);
and AND3 (N489, N485, N16, N106);
not NOT1 (N490, N489);
buf BUF1 (N491, N484);
xor XOR2 (N492, N486, N72);
not NOT1 (N493, N490);
or OR2 (N494, N477, N81);
nor NOR4 (N495, N492, N347, N23, N145);
xor XOR2 (N496, N494, N168);
buf BUF1 (N497, N496);
not NOT1 (N498, N482);
buf BUF1 (N499, N491);
or OR2 (N500, N499, N326);
and AND2 (N501, N497, N355);
not NOT1 (N502, N501);
nand NAND2 (N503, N488, N445);
xor XOR2 (N504, N480, N389);
nand NAND3 (N505, N487, N275, N73);
xor XOR2 (N506, N495, N17);
nand NAND4 (N507, N475, N144, N308, N172);
not NOT1 (N508, N505);
not NOT1 (N509, N508);
not NOT1 (N510, N503);
buf BUF1 (N511, N509);
buf BUF1 (N512, N511);
xor XOR2 (N513, N500, N236);
nor NOR3 (N514, N493, N207, N345);
and AND3 (N515, N513, N177, N384);
nor NOR3 (N516, N504, N163, N242);
nand NAND4 (N517, N507, N26, N328, N294);
nand NAND3 (N518, N502, N260, N150);
and AND3 (N519, N483, N14, N30);
endmodule