// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23;

output N16017,N16022,N16013,N16015,N16003,N16019,N16011,N15993,N16021,N16023;

not NOT1 (N24, N7);
not NOT1 (N25, N17);
or OR2 (N26, N10, N13);
or OR2 (N27, N16, N4);
buf BUF1 (N28, N12);
buf BUF1 (N29, N11);
xor XOR2 (N30, N29, N14);
and AND4 (N31, N8, N24, N24, N13);
not NOT1 (N32, N24);
xor XOR2 (N33, N4, N29);
buf BUF1 (N34, N18);
not NOT1 (N35, N9);
nand NAND3 (N36, N26, N32, N23);
not NOT1 (N37, N29);
nand NAND2 (N38, N35, N6);
buf BUF1 (N39, N34);
not NOT1 (N40, N39);
or OR2 (N41, N33, N10);
buf BUF1 (N42, N31);
nand NAND2 (N43, N40, N8);
nand NAND4 (N44, N41, N43, N16, N23);
or OR4 (N45, N43, N43, N24, N41);
nor NOR2 (N46, N30, N37);
nand NAND2 (N47, N43, N2);
not NOT1 (N48, N45);
not NOT1 (N49, N27);
or OR4 (N50, N38, N43, N10, N16);
and AND4 (N51, N25, N7, N19, N15);
or OR3 (N52, N36, N21, N17);
nand NAND4 (N53, N42, N4, N16, N44);
buf BUF1 (N54, N15);
buf BUF1 (N55, N47);
and AND4 (N56, N48, N43, N43, N48);
buf BUF1 (N57, N46);
xor XOR2 (N58, N49, N18);
not NOT1 (N59, N54);
buf BUF1 (N60, N56);
or OR4 (N61, N57, N29, N27, N35);
nor NOR3 (N62, N58, N7, N47);
nor NOR4 (N63, N53, N43, N6, N54);
and AND4 (N64, N62, N34, N53, N33);
not NOT1 (N65, N52);
nor NOR2 (N66, N60, N63);
not NOT1 (N67, N61);
and AND4 (N68, N58, N20, N64, N8);
nand NAND2 (N69, N37, N31);
nand NAND3 (N70, N59, N69, N26);
or OR4 (N71, N45, N43, N51, N49);
or OR4 (N72, N41, N32, N52, N8);
nor NOR3 (N73, N68, N31, N18);
or OR3 (N74, N50, N46, N40);
not NOT1 (N75, N74);
and AND3 (N76, N73, N36, N31);
and AND4 (N77, N66, N36, N45, N8);
not NOT1 (N78, N76);
xor XOR2 (N79, N78, N36);
xor XOR2 (N80, N55, N9);
and AND4 (N81, N71, N15, N4, N31);
buf BUF1 (N82, N72);
or OR2 (N83, N80, N69);
and AND4 (N84, N28, N70, N49, N37);
and AND3 (N85, N20, N39, N38);
or OR2 (N86, N81, N7);
and AND3 (N87, N82, N83, N49);
buf BUF1 (N88, N22);
xor XOR2 (N89, N75, N76);
and AND4 (N90, N65, N42, N59, N13);
buf BUF1 (N91, N79);
not NOT1 (N92, N86);
and AND4 (N93, N91, N15, N1, N12);
buf BUF1 (N94, N67);
buf BUF1 (N95, N88);
nand NAND3 (N96, N94, N27, N78);
nand NAND3 (N97, N92, N23, N42);
or OR4 (N98, N90, N30, N1, N70);
buf BUF1 (N99, N87);
xor XOR2 (N100, N97, N9);
or OR4 (N101, N85, N30, N22, N52);
nand NAND2 (N102, N89, N77);
and AND2 (N103, N93, N16);
buf BUF1 (N104, N34);
not NOT1 (N105, N98);
and AND3 (N106, N95, N89, N20);
nand NAND3 (N107, N104, N90, N24);
and AND2 (N108, N101, N16);
nand NAND4 (N109, N103, N10, N106, N65);
and AND2 (N110, N104, N91);
xor XOR2 (N111, N108, N6);
nand NAND2 (N112, N111, N2);
or OR2 (N113, N102, N72);
not NOT1 (N114, N110);
xor XOR2 (N115, N112, N35);
buf BUF1 (N116, N115);
not NOT1 (N117, N107);
nor NOR3 (N118, N84, N74, N8);
and AND4 (N119, N117, N83, N36, N48);
nor NOR2 (N120, N96, N85);
nand NAND4 (N121, N114, N96, N110, N40);
nor NOR4 (N122, N116, N13, N65, N40);
nor NOR4 (N123, N121, N101, N28, N7);
nor NOR4 (N124, N113, N117, N47, N31);
not NOT1 (N125, N124);
not NOT1 (N126, N122);
or OR3 (N127, N105, N124, N10);
xor XOR2 (N128, N123, N15);
nand NAND4 (N129, N100, N83, N70, N62);
not NOT1 (N130, N99);
not NOT1 (N131, N130);
and AND2 (N132, N120, N106);
and AND3 (N133, N126, N38, N61);
buf BUF1 (N134, N125);
buf BUF1 (N135, N132);
not NOT1 (N136, N128);
nand NAND3 (N137, N134, N134, N131);
not NOT1 (N138, N118);
nand NAND4 (N139, N4, N34, N89, N1);
nor NOR3 (N140, N127, N82, N53);
and AND3 (N141, N133, N60, N86);
and AND4 (N142, N119, N93, N114, N141);
nor NOR2 (N143, N112, N16);
buf BUF1 (N144, N143);
nand NAND4 (N145, N140, N42, N32, N110);
buf BUF1 (N146, N137);
nor NOR2 (N147, N136, N48);
nand NAND2 (N148, N129, N46);
nand NAND3 (N149, N139, N18, N118);
or OR2 (N150, N138, N20);
nor NOR4 (N151, N147, N98, N104, N39);
nand NAND4 (N152, N146, N80, N136, N141);
xor XOR2 (N153, N149, N24);
or OR4 (N154, N151, N32, N109, N72);
nor NOR3 (N155, N10, N64, N21);
and AND4 (N156, N155, N72, N1, N130);
nand NAND3 (N157, N145, N83, N23);
nand NAND3 (N158, N152, N42, N18);
nor NOR3 (N159, N157, N25, N70);
xor XOR2 (N160, N158, N1);
or OR4 (N161, N144, N23, N139, N111);
nand NAND2 (N162, N153, N11);
xor XOR2 (N163, N135, N145);
not NOT1 (N164, N159);
and AND4 (N165, N160, N91, N148, N144);
or OR4 (N166, N53, N99, N123, N45);
buf BUF1 (N167, N161);
nor NOR3 (N168, N142, N90, N123);
and AND2 (N169, N166, N131);
not NOT1 (N170, N150);
and AND2 (N171, N164, N50);
and AND4 (N172, N167, N75, N1, N123);
and AND3 (N173, N168, N86, N161);
or OR3 (N174, N162, N106, N5);
or OR2 (N175, N173, N50);
nor NOR4 (N176, N170, N55, N75, N21);
buf BUF1 (N177, N174);
not NOT1 (N178, N172);
not NOT1 (N179, N163);
nor NOR2 (N180, N179, N60);
and AND3 (N181, N177, N159, N124);
xor XOR2 (N182, N176, N24);
xor XOR2 (N183, N171, N34);
xor XOR2 (N184, N165, N73);
xor XOR2 (N185, N156, N69);
xor XOR2 (N186, N185, N81);
not NOT1 (N187, N182);
nor NOR4 (N188, N183, N94, N162, N47);
and AND2 (N189, N180, N54);
not NOT1 (N190, N187);
buf BUF1 (N191, N181);
nor NOR2 (N192, N189, N87);
nand NAND3 (N193, N192, N110, N33);
buf BUF1 (N194, N154);
nand NAND3 (N195, N186, N120, N90);
nor NOR3 (N196, N194, N25, N24);
or OR4 (N197, N169, N158, N21, N4);
nand NAND2 (N198, N195, N94);
nand NAND2 (N199, N197, N150);
not NOT1 (N200, N196);
nand NAND3 (N201, N191, N35, N92);
nand NAND3 (N202, N199, N121, N116);
not NOT1 (N203, N193);
nand NAND4 (N204, N190, N3, N130, N185);
nand NAND4 (N205, N201, N164, N171, N48);
and AND4 (N206, N188, N8, N192, N96);
xor XOR2 (N207, N203, N148);
buf BUF1 (N208, N200);
and AND2 (N209, N178, N164);
nor NOR3 (N210, N209, N121, N186);
or OR4 (N211, N205, N36, N88, N26);
nand NAND4 (N212, N202, N143, N187, N184);
xor XOR2 (N213, N151, N211);
buf BUF1 (N214, N81);
and AND3 (N215, N206, N127, N97);
xor XOR2 (N216, N207, N190);
not NOT1 (N217, N216);
nor NOR2 (N218, N213, N169);
not NOT1 (N219, N217);
or OR2 (N220, N215, N167);
nor NOR3 (N221, N198, N138, N95);
buf BUF1 (N222, N204);
buf BUF1 (N223, N218);
and AND4 (N224, N208, N129, N56, N35);
xor XOR2 (N225, N210, N105);
xor XOR2 (N226, N222, N217);
and AND2 (N227, N212, N23);
and AND3 (N228, N221, N9, N190);
and AND4 (N229, N225, N101, N50, N92);
buf BUF1 (N230, N214);
and AND4 (N231, N219, N180, N212, N85);
not NOT1 (N232, N227);
buf BUF1 (N233, N228);
nor NOR3 (N234, N175, N28, N155);
not NOT1 (N235, N231);
and AND2 (N236, N233, N19);
and AND3 (N237, N235, N57, N201);
buf BUF1 (N238, N237);
nand NAND2 (N239, N236, N199);
or OR2 (N240, N226, N216);
or OR2 (N241, N230, N153);
buf BUF1 (N242, N224);
buf BUF1 (N243, N232);
xor XOR2 (N244, N229, N171);
buf BUF1 (N245, N243);
or OR4 (N246, N238, N238, N13, N140);
or OR3 (N247, N240, N228, N69);
nand NAND2 (N248, N244, N105);
nor NOR4 (N249, N241, N108, N245, N149);
not NOT1 (N250, N209);
nand NAND2 (N251, N234, N61);
nor NOR4 (N252, N250, N151, N11, N30);
and AND3 (N253, N249, N156, N127);
or OR3 (N254, N220, N158, N45);
nor NOR2 (N255, N239, N19);
nor NOR3 (N256, N254, N99, N204);
nor NOR4 (N257, N256, N127, N135, N42);
nand NAND3 (N258, N242, N186, N208);
nand NAND2 (N259, N248, N14);
not NOT1 (N260, N259);
buf BUF1 (N261, N258);
or OR4 (N262, N223, N31, N178, N72);
nor NOR4 (N263, N260, N39, N25, N23);
nor NOR4 (N264, N251, N198, N28, N172);
nor NOR3 (N265, N262, N250, N139);
buf BUF1 (N266, N264);
and AND4 (N267, N266, N230, N213, N135);
not NOT1 (N268, N261);
nand NAND2 (N269, N247, N266);
not NOT1 (N270, N263);
or OR3 (N271, N268, N234, N248);
buf BUF1 (N272, N267);
xor XOR2 (N273, N272, N270);
not NOT1 (N274, N206);
nand NAND4 (N275, N252, N90, N195, N169);
or OR3 (N276, N271, N9, N90);
not NOT1 (N277, N273);
nand NAND2 (N278, N277, N204);
not NOT1 (N279, N269);
and AND2 (N280, N276, N62);
and AND2 (N281, N246, N125);
and AND2 (N282, N280, N259);
buf BUF1 (N283, N257);
buf BUF1 (N284, N281);
xor XOR2 (N285, N274, N266);
or OR2 (N286, N279, N12);
buf BUF1 (N287, N286);
buf BUF1 (N288, N282);
xor XOR2 (N289, N265, N147);
nand NAND2 (N290, N289, N253);
buf BUF1 (N291, N134);
or OR2 (N292, N284, N37);
and AND3 (N293, N275, N260, N159);
or OR2 (N294, N290, N291);
nand NAND3 (N295, N3, N42, N121);
and AND3 (N296, N278, N32, N101);
buf BUF1 (N297, N285);
nor NOR4 (N298, N288, N116, N96, N288);
not NOT1 (N299, N296);
not NOT1 (N300, N297);
or OR2 (N301, N298, N10);
xor XOR2 (N302, N255, N110);
xor XOR2 (N303, N299, N61);
xor XOR2 (N304, N293, N224);
or OR2 (N305, N301, N134);
nand NAND4 (N306, N295, N241, N67, N182);
not NOT1 (N307, N305);
not NOT1 (N308, N292);
and AND3 (N309, N306, N239, N183);
xor XOR2 (N310, N287, N180);
nor NOR4 (N311, N308, N36, N240, N244);
not NOT1 (N312, N283);
nor NOR3 (N313, N303, N244, N217);
buf BUF1 (N314, N311);
xor XOR2 (N315, N304, N216);
nor NOR3 (N316, N314, N157, N220);
buf BUF1 (N317, N316);
and AND2 (N318, N317, N208);
buf BUF1 (N319, N313);
xor XOR2 (N320, N318, N141);
or OR4 (N321, N312, N129, N111, N169);
nor NOR2 (N322, N300, N1);
nor NOR2 (N323, N315, N131);
and AND4 (N324, N310, N241, N228, N240);
not NOT1 (N325, N302);
not NOT1 (N326, N309);
and AND3 (N327, N322, N240, N267);
nand NAND2 (N328, N323, N266);
nor NOR3 (N329, N327, N218, N9);
or OR4 (N330, N326, N168, N137, N141);
xor XOR2 (N331, N329, N77);
and AND4 (N332, N325, N191, N239, N251);
buf BUF1 (N333, N332);
not NOT1 (N334, N330);
xor XOR2 (N335, N319, N319);
nand NAND4 (N336, N333, N185, N307, N130);
or OR3 (N337, N267, N165, N152);
buf BUF1 (N338, N335);
and AND4 (N339, N337, N24, N202, N180);
and AND3 (N340, N334, N232, N338);
nand NAND3 (N341, N206, N177, N299);
xor XOR2 (N342, N341, N126);
and AND3 (N343, N331, N60, N117);
buf BUF1 (N344, N324);
nor NOR2 (N345, N320, N22);
nand NAND3 (N346, N345, N44, N246);
and AND2 (N347, N294, N87);
and AND2 (N348, N344, N24);
buf BUF1 (N349, N328);
buf BUF1 (N350, N340);
nand NAND3 (N351, N348, N147, N228);
nor NOR4 (N352, N351, N253, N291, N55);
not NOT1 (N353, N350);
and AND4 (N354, N352, N351, N6, N224);
nor NOR4 (N355, N342, N284, N258, N270);
or OR3 (N356, N354, N213, N339);
not NOT1 (N357, N344);
buf BUF1 (N358, N356);
nor NOR3 (N359, N358, N153, N262);
xor XOR2 (N360, N353, N22);
nor NOR2 (N361, N347, N50);
not NOT1 (N362, N361);
and AND4 (N363, N321, N42, N262, N155);
or OR4 (N364, N349, N17, N353, N31);
xor XOR2 (N365, N363, N126);
buf BUF1 (N366, N336);
nand NAND4 (N367, N364, N266, N125, N327);
xor XOR2 (N368, N346, N132);
xor XOR2 (N369, N365, N255);
not NOT1 (N370, N367);
nor NOR4 (N371, N370, N129, N282, N306);
nand NAND4 (N372, N355, N261, N175, N70);
nand NAND4 (N373, N357, N251, N151, N152);
not NOT1 (N374, N362);
or OR3 (N375, N360, N1, N279);
nand NAND2 (N376, N359, N320);
nand NAND2 (N377, N371, N19);
not NOT1 (N378, N374);
nand NAND2 (N379, N375, N120);
or OR3 (N380, N373, N318, N280);
xor XOR2 (N381, N366, N329);
or OR2 (N382, N377, N207);
nand NAND3 (N383, N343, N170, N42);
xor XOR2 (N384, N376, N283);
xor XOR2 (N385, N379, N151);
nor NOR3 (N386, N381, N300, N53);
buf BUF1 (N387, N383);
not NOT1 (N388, N387);
and AND3 (N389, N386, N275, N248);
or OR2 (N390, N389, N385);
buf BUF1 (N391, N317);
and AND4 (N392, N368, N300, N143, N165);
xor XOR2 (N393, N390, N58);
nor NOR2 (N394, N392, N308);
and AND3 (N395, N394, N116, N353);
buf BUF1 (N396, N391);
not NOT1 (N397, N372);
nand NAND4 (N398, N396, N70, N198, N351);
not NOT1 (N399, N395);
buf BUF1 (N400, N399);
xor XOR2 (N401, N382, N29);
nor NOR2 (N402, N400, N350);
buf BUF1 (N403, N369);
or OR2 (N404, N378, N185);
xor XOR2 (N405, N388, N355);
not NOT1 (N406, N397);
not NOT1 (N407, N406);
not NOT1 (N408, N380);
not NOT1 (N409, N398);
nand NAND4 (N410, N393, N175, N201, N409);
xor XOR2 (N411, N4, N185);
nor NOR3 (N412, N404, N311, N220);
or OR4 (N413, N384, N274, N112, N70);
buf BUF1 (N414, N407);
xor XOR2 (N415, N412, N28);
or OR2 (N416, N413, N359);
nand NAND4 (N417, N405, N247, N262, N374);
nand NAND4 (N418, N411, N233, N297, N56);
nand NAND2 (N419, N414, N371);
or OR4 (N420, N403, N302, N167, N291);
nor NOR4 (N421, N416, N8, N351, N237);
and AND2 (N422, N417, N133);
nor NOR3 (N423, N415, N185, N174);
not NOT1 (N424, N401);
nor NOR3 (N425, N420, N376, N359);
or OR4 (N426, N422, N315, N346, N209);
and AND4 (N427, N410, N191, N47, N392);
not NOT1 (N428, N423);
nand NAND4 (N429, N426, N67, N212, N141);
buf BUF1 (N430, N419);
and AND2 (N431, N427, N166);
and AND4 (N432, N428, N13, N41, N272);
nand NAND2 (N433, N421, N261);
nor NOR3 (N434, N424, N196, N185);
buf BUF1 (N435, N431);
or OR3 (N436, N430, N6, N273);
not NOT1 (N437, N434);
nand NAND2 (N438, N418, N137);
or OR2 (N439, N425, N165);
and AND3 (N440, N439, N295, N200);
nand NAND2 (N441, N408, N32);
buf BUF1 (N442, N437);
nand NAND2 (N443, N429, N140);
buf BUF1 (N444, N435);
nor NOR3 (N445, N402, N371, N243);
nand NAND2 (N446, N438, N60);
nand NAND3 (N447, N443, N50, N354);
or OR4 (N448, N432, N172, N18, N156);
nand NAND4 (N449, N448, N318, N225, N431);
nor NOR3 (N450, N447, N211, N19);
not NOT1 (N451, N440);
or OR3 (N452, N450, N162, N417);
not NOT1 (N453, N444);
xor XOR2 (N454, N436, N209);
nand NAND2 (N455, N441, N237);
buf BUF1 (N456, N451);
nor NOR3 (N457, N433, N23, N407);
or OR4 (N458, N449, N279, N146, N341);
xor XOR2 (N459, N453, N253);
buf BUF1 (N460, N456);
xor XOR2 (N461, N459, N194);
xor XOR2 (N462, N445, N134);
xor XOR2 (N463, N458, N201);
not NOT1 (N464, N457);
and AND2 (N465, N446, N12);
or OR3 (N466, N462, N1, N123);
or OR3 (N467, N465, N291, N263);
xor XOR2 (N468, N463, N295);
buf BUF1 (N469, N460);
and AND2 (N470, N468, N270);
nor NOR3 (N471, N467, N101, N252);
buf BUF1 (N472, N454);
and AND4 (N473, N464, N344, N60, N294);
xor XOR2 (N474, N452, N376);
nor NOR2 (N475, N469, N370);
nor NOR4 (N476, N471, N177, N441, N196);
and AND3 (N477, N474, N467, N340);
nor NOR4 (N478, N470, N82, N63, N342);
nand NAND4 (N479, N473, N30, N188, N441);
buf BUF1 (N480, N461);
not NOT1 (N481, N442);
xor XOR2 (N482, N466, N431);
buf BUF1 (N483, N479);
or OR4 (N484, N480, N448, N284, N300);
not NOT1 (N485, N478);
buf BUF1 (N486, N475);
xor XOR2 (N487, N482, N287);
buf BUF1 (N488, N486);
and AND3 (N489, N477, N308, N68);
not NOT1 (N490, N485);
or OR2 (N491, N476, N398);
or OR2 (N492, N489, N28);
nor NOR3 (N493, N481, N446, N386);
nor NOR2 (N494, N492, N409);
xor XOR2 (N495, N472, N56);
or OR2 (N496, N455, N125);
nor NOR2 (N497, N496, N66);
not NOT1 (N498, N488);
and AND4 (N499, N497, N291, N234, N432);
nor NOR3 (N500, N495, N151, N356);
nand NAND4 (N501, N498, N494, N106, N16);
or OR4 (N502, N394, N23, N160, N20);
buf BUF1 (N503, N502);
nor NOR4 (N504, N491, N294, N254, N108);
or OR2 (N505, N503, N108);
xor XOR2 (N506, N505, N383);
buf BUF1 (N507, N483);
nor NOR4 (N508, N501, N447, N325, N33);
nor NOR2 (N509, N504, N18);
and AND4 (N510, N508, N12, N113, N418);
buf BUF1 (N511, N507);
or OR4 (N512, N510, N96, N422, N263);
not NOT1 (N513, N490);
nand NAND3 (N514, N511, N387, N369);
xor XOR2 (N515, N487, N198);
xor XOR2 (N516, N513, N296);
xor XOR2 (N517, N515, N116);
nand NAND3 (N518, N506, N423, N322);
or OR2 (N519, N512, N295);
nor NOR4 (N520, N518, N209, N514, N67);
xor XOR2 (N521, N467, N127);
nor NOR3 (N522, N493, N19, N448);
not NOT1 (N523, N500);
buf BUF1 (N524, N519);
not NOT1 (N525, N520);
or OR2 (N526, N484, N179);
or OR4 (N527, N521, N3, N15, N89);
nand NAND4 (N528, N516, N468, N260, N279);
nand NAND4 (N529, N509, N289, N506, N89);
xor XOR2 (N530, N528, N451);
xor XOR2 (N531, N499, N380);
not NOT1 (N532, N526);
nor NOR3 (N533, N530, N507, N3);
not NOT1 (N534, N531);
and AND4 (N535, N532, N479, N399, N261);
xor XOR2 (N536, N534, N218);
buf BUF1 (N537, N523);
and AND4 (N538, N537, N536, N276, N359);
or OR2 (N539, N48, N419);
not NOT1 (N540, N539);
or OR2 (N541, N538, N144);
not NOT1 (N542, N522);
nor NOR4 (N543, N524, N446, N470, N397);
nor NOR4 (N544, N543, N384, N58, N144);
not NOT1 (N545, N541);
nand NAND2 (N546, N529, N378);
and AND3 (N547, N540, N377, N524);
or OR4 (N548, N547, N424, N436, N364);
nor NOR2 (N549, N527, N38);
not NOT1 (N550, N525);
not NOT1 (N551, N550);
nand NAND4 (N552, N517, N156, N2, N338);
and AND3 (N553, N533, N311, N111);
nand NAND2 (N554, N545, N8);
or OR4 (N555, N552, N109, N354, N272);
xor XOR2 (N556, N535, N452);
xor XOR2 (N557, N554, N290);
not NOT1 (N558, N553);
nor NOR3 (N559, N544, N531, N56);
and AND4 (N560, N559, N478, N141, N347);
nand NAND3 (N561, N556, N101, N536);
nand NAND2 (N562, N555, N58);
not NOT1 (N563, N549);
nand NAND2 (N564, N542, N317);
nor NOR2 (N565, N563, N409);
nand NAND3 (N566, N546, N125, N64);
nor NOR3 (N567, N561, N393, N537);
xor XOR2 (N568, N548, N373);
not NOT1 (N569, N560);
or OR2 (N570, N564, N312);
nand NAND4 (N571, N566, N324, N428, N167);
not NOT1 (N572, N557);
or OR3 (N573, N567, N421, N481);
nand NAND4 (N574, N568, N217, N263, N408);
and AND2 (N575, N565, N367);
xor XOR2 (N576, N575, N185);
nor NOR2 (N577, N572, N113);
or OR2 (N578, N576, N145);
nand NAND3 (N579, N562, N309, N568);
xor XOR2 (N580, N578, N28);
buf BUF1 (N581, N573);
buf BUF1 (N582, N581);
buf BUF1 (N583, N582);
buf BUF1 (N584, N569);
and AND3 (N585, N574, N407, N475);
nand NAND4 (N586, N571, N532, N549, N449);
nand NAND2 (N587, N584, N580);
not NOT1 (N588, N245);
and AND4 (N589, N587, N377, N197, N493);
xor XOR2 (N590, N585, N244);
not NOT1 (N591, N586);
not NOT1 (N592, N558);
nand NAND2 (N593, N577, N282);
nor NOR4 (N594, N591, N387, N363, N214);
nand NAND3 (N595, N590, N77, N512);
nor NOR2 (N596, N594, N427);
or OR3 (N597, N589, N172, N432);
xor XOR2 (N598, N595, N592);
nor NOR4 (N599, N436, N451, N128, N392);
nand NAND2 (N600, N599, N57);
not NOT1 (N601, N551);
and AND2 (N602, N601, N247);
xor XOR2 (N603, N598, N206);
nand NAND4 (N604, N579, N459, N489, N85);
nand NAND2 (N605, N602, N415);
buf BUF1 (N606, N600);
xor XOR2 (N607, N570, N513);
nand NAND2 (N608, N605, N161);
and AND2 (N609, N603, N458);
and AND4 (N610, N596, N139, N223, N504);
or OR3 (N611, N597, N581, N493);
nor NOR2 (N612, N583, N529);
and AND2 (N613, N611, N481);
not NOT1 (N614, N588);
and AND3 (N615, N609, N265, N612);
nor NOR4 (N616, N305, N478, N113, N402);
nand NAND2 (N617, N613, N469);
nand NAND3 (N618, N593, N590, N320);
buf BUF1 (N619, N615);
nor NOR4 (N620, N616, N356, N185, N170);
not NOT1 (N621, N619);
nand NAND2 (N622, N607, N361);
xor XOR2 (N623, N610, N111);
nor NOR4 (N624, N606, N569, N556, N99);
or OR3 (N625, N620, N311, N416);
xor XOR2 (N626, N614, N22);
not NOT1 (N627, N624);
nand NAND2 (N628, N625, N129);
nor NOR2 (N629, N618, N413);
buf BUF1 (N630, N622);
nand NAND3 (N631, N626, N289, N431);
and AND2 (N632, N627, N351);
buf BUF1 (N633, N621);
not NOT1 (N634, N632);
nor NOR4 (N635, N604, N381, N345, N156);
nand NAND2 (N636, N629, N471);
and AND4 (N637, N631, N528, N384, N466);
buf BUF1 (N638, N636);
buf BUF1 (N639, N628);
nor NOR3 (N640, N630, N229, N171);
not NOT1 (N641, N635);
nor NOR4 (N642, N623, N32, N368, N123);
not NOT1 (N643, N641);
nand NAND2 (N644, N639, N405);
buf BUF1 (N645, N638);
or OR4 (N646, N645, N645, N315, N81);
xor XOR2 (N647, N640, N201);
nor NOR3 (N648, N634, N518, N385);
buf BUF1 (N649, N643);
not NOT1 (N650, N633);
xor XOR2 (N651, N648, N127);
nand NAND4 (N652, N646, N551, N414, N219);
and AND4 (N653, N647, N252, N396, N164);
or OR2 (N654, N642, N578);
nand NAND4 (N655, N653, N111, N324, N417);
not NOT1 (N656, N649);
buf BUF1 (N657, N656);
nand NAND3 (N658, N657, N175, N636);
not NOT1 (N659, N655);
buf BUF1 (N660, N658);
not NOT1 (N661, N650);
nand NAND2 (N662, N659, N435);
nand NAND3 (N663, N617, N592, N112);
nor NOR2 (N664, N644, N454);
and AND2 (N665, N608, N262);
nand NAND4 (N666, N663, N302, N39, N283);
nor NOR4 (N667, N666, N570, N130, N218);
nand NAND3 (N668, N667, N381, N495);
nor NOR3 (N669, N654, N279, N527);
and AND4 (N670, N664, N341, N256, N615);
nand NAND2 (N671, N651, N425);
nand NAND2 (N672, N661, N396);
or OR4 (N673, N652, N392, N1, N477);
xor XOR2 (N674, N672, N307);
not NOT1 (N675, N669);
buf BUF1 (N676, N637);
or OR3 (N677, N675, N101, N285);
xor XOR2 (N678, N674, N21);
xor XOR2 (N679, N678, N117);
buf BUF1 (N680, N670);
nand NAND3 (N681, N665, N327, N364);
not NOT1 (N682, N668);
or OR2 (N683, N676, N394);
nor NOR4 (N684, N671, N337, N164, N122);
buf BUF1 (N685, N679);
not NOT1 (N686, N682);
nor NOR3 (N687, N677, N630, N193);
xor XOR2 (N688, N684, N162);
not NOT1 (N689, N680);
nor NOR4 (N690, N660, N231, N211, N383);
xor XOR2 (N691, N686, N214);
nand NAND3 (N692, N662, N69, N542);
buf BUF1 (N693, N690);
xor XOR2 (N694, N685, N262);
buf BUF1 (N695, N691);
nor NOR4 (N696, N687, N509, N569, N143);
nand NAND2 (N697, N673, N13);
buf BUF1 (N698, N692);
nand NAND4 (N699, N695, N476, N122, N577);
and AND4 (N700, N689, N79, N521, N393);
nor NOR2 (N701, N696, N544);
xor XOR2 (N702, N681, N54);
buf BUF1 (N703, N688);
buf BUF1 (N704, N697);
nand NAND2 (N705, N700, N124);
not NOT1 (N706, N693);
nor NOR3 (N707, N705, N568, N324);
buf BUF1 (N708, N707);
and AND3 (N709, N708, N249, N672);
or OR3 (N710, N701, N60, N334);
and AND4 (N711, N703, N247, N240, N483);
and AND2 (N712, N683, N692);
nor NOR4 (N713, N699, N87, N243, N361);
nor NOR3 (N714, N702, N68, N705);
or OR2 (N715, N706, N59);
and AND3 (N716, N698, N576, N3);
or OR3 (N717, N709, N480, N670);
and AND2 (N718, N712, N108);
or OR2 (N719, N718, N174);
xor XOR2 (N720, N694, N359);
and AND3 (N721, N711, N283, N292);
nand NAND3 (N722, N719, N186, N430);
nand NAND2 (N723, N721, N481);
not NOT1 (N724, N717);
nor NOR4 (N725, N723, N286, N348, N77);
and AND3 (N726, N725, N9, N138);
nand NAND3 (N727, N720, N286, N82);
or OR2 (N728, N710, N686);
or OR2 (N729, N713, N579);
xor XOR2 (N730, N722, N62);
and AND2 (N731, N728, N149);
buf BUF1 (N732, N704);
and AND3 (N733, N715, N154, N361);
xor XOR2 (N734, N730, N626);
xor XOR2 (N735, N731, N542);
buf BUF1 (N736, N735);
and AND2 (N737, N736, N373);
buf BUF1 (N738, N733);
buf BUF1 (N739, N727);
or OR2 (N740, N716, N289);
and AND2 (N741, N737, N585);
not NOT1 (N742, N729);
nand NAND3 (N743, N738, N13, N389);
or OR2 (N744, N741, N573);
buf BUF1 (N745, N743);
and AND4 (N746, N739, N633, N96, N737);
xor XOR2 (N747, N724, N170);
nor NOR3 (N748, N745, N549, N657);
not NOT1 (N749, N742);
not NOT1 (N750, N732);
buf BUF1 (N751, N740);
nand NAND4 (N752, N747, N34, N319, N207);
xor XOR2 (N753, N750, N623);
xor XOR2 (N754, N752, N505);
or OR3 (N755, N714, N16, N585);
and AND4 (N756, N754, N546, N16, N686);
not NOT1 (N757, N749);
buf BUF1 (N758, N755);
buf BUF1 (N759, N753);
nor NOR3 (N760, N734, N451, N432);
buf BUF1 (N761, N758);
and AND3 (N762, N726, N613, N319);
nor NOR2 (N763, N756, N603);
not NOT1 (N764, N748);
nand NAND2 (N765, N759, N492);
buf BUF1 (N766, N763);
or OR4 (N767, N757, N288, N760, N471);
and AND2 (N768, N574, N581);
buf BUF1 (N769, N761);
xor XOR2 (N770, N766, N458);
xor XOR2 (N771, N746, N154);
nor NOR3 (N772, N744, N111, N190);
nor NOR3 (N773, N769, N732, N620);
xor XOR2 (N774, N762, N6);
and AND3 (N775, N770, N165, N120);
or OR4 (N776, N772, N575, N304, N125);
xor XOR2 (N777, N751, N301);
xor XOR2 (N778, N771, N624);
xor XOR2 (N779, N778, N510);
nor NOR2 (N780, N779, N314);
or OR4 (N781, N777, N743, N432, N410);
xor XOR2 (N782, N781, N259);
not NOT1 (N783, N780);
or OR4 (N784, N767, N361, N2, N72);
or OR3 (N785, N768, N706, N448);
xor XOR2 (N786, N784, N150);
xor XOR2 (N787, N782, N472);
not NOT1 (N788, N774);
nor NOR2 (N789, N764, N646);
buf BUF1 (N790, N776);
or OR4 (N791, N773, N283, N643, N182);
and AND4 (N792, N787, N8, N94, N598);
nand NAND2 (N793, N783, N322);
not NOT1 (N794, N791);
and AND3 (N795, N792, N410, N558);
not NOT1 (N796, N786);
not NOT1 (N797, N785);
xor XOR2 (N798, N765, N573);
nand NAND4 (N799, N789, N298, N608, N48);
not NOT1 (N800, N795);
and AND3 (N801, N788, N417, N761);
xor XOR2 (N802, N797, N426);
buf BUF1 (N803, N775);
buf BUF1 (N804, N793);
nor NOR4 (N805, N801, N334, N6, N775);
nand NAND4 (N806, N800, N169, N606, N279);
xor XOR2 (N807, N790, N455);
nand NAND4 (N808, N804, N297, N725, N232);
and AND4 (N809, N802, N501, N197, N787);
or OR3 (N810, N796, N528, N561);
not NOT1 (N811, N799);
buf BUF1 (N812, N794);
or OR4 (N813, N806, N462, N635, N439);
nor NOR2 (N814, N807, N317);
nor NOR2 (N815, N803, N184);
nor NOR4 (N816, N798, N571, N317, N684);
nand NAND2 (N817, N805, N43);
not NOT1 (N818, N815);
nand NAND2 (N819, N808, N237);
and AND3 (N820, N812, N814, N783);
not NOT1 (N821, N591);
nor NOR2 (N822, N817, N78);
not NOT1 (N823, N820);
and AND3 (N824, N822, N372, N313);
not NOT1 (N825, N811);
not NOT1 (N826, N810);
and AND3 (N827, N819, N693, N314);
and AND4 (N828, N823, N769, N32, N494);
and AND4 (N829, N816, N178, N647, N613);
and AND3 (N830, N828, N532, N416);
buf BUF1 (N831, N827);
and AND3 (N832, N825, N55, N40);
nor NOR4 (N833, N830, N193, N203, N49);
not NOT1 (N834, N833);
not NOT1 (N835, N818);
buf BUF1 (N836, N826);
and AND2 (N837, N836, N67);
xor XOR2 (N838, N824, N378);
not NOT1 (N839, N835);
nor NOR2 (N840, N813, N340);
nor NOR3 (N841, N840, N761, N210);
or OR2 (N842, N837, N623);
not NOT1 (N843, N834);
and AND4 (N844, N841, N700, N536, N221);
xor XOR2 (N845, N842, N622);
xor XOR2 (N846, N845, N443);
nand NAND2 (N847, N809, N402);
buf BUF1 (N848, N839);
and AND3 (N849, N846, N19, N777);
buf BUF1 (N850, N844);
or OR2 (N851, N849, N509);
nor NOR3 (N852, N847, N334, N676);
buf BUF1 (N853, N832);
xor XOR2 (N854, N852, N459);
buf BUF1 (N855, N843);
nand NAND2 (N856, N850, N492);
buf BUF1 (N857, N855);
nor NOR3 (N858, N829, N854, N678);
and AND3 (N859, N711, N853, N440);
nand NAND4 (N860, N667, N606, N24, N205);
and AND4 (N861, N859, N247, N723, N462);
xor XOR2 (N862, N821, N685);
nor NOR3 (N863, N862, N410, N777);
not NOT1 (N864, N856);
nor NOR2 (N865, N831, N840);
not NOT1 (N866, N861);
buf BUF1 (N867, N866);
nand NAND3 (N868, N860, N218, N209);
nor NOR2 (N869, N857, N96);
not NOT1 (N870, N848);
nand NAND3 (N871, N864, N204, N360);
buf BUF1 (N872, N858);
or OR4 (N873, N838, N268, N613, N263);
or OR3 (N874, N871, N577, N18);
xor XOR2 (N875, N865, N566);
xor XOR2 (N876, N851, N80);
nor NOR2 (N877, N870, N364);
nor NOR2 (N878, N872, N60);
nor NOR2 (N879, N873, N117);
not NOT1 (N880, N877);
buf BUF1 (N881, N878);
or OR3 (N882, N868, N514, N795);
nand NAND2 (N883, N869, N870);
nor NOR3 (N884, N876, N14, N687);
not NOT1 (N885, N874);
or OR2 (N886, N863, N872);
xor XOR2 (N887, N879, N260);
nand NAND2 (N888, N883, N565);
nand NAND4 (N889, N887, N802, N647, N216);
not NOT1 (N890, N886);
buf BUF1 (N891, N882);
or OR2 (N892, N875, N768);
not NOT1 (N893, N884);
xor XOR2 (N894, N888, N878);
buf BUF1 (N895, N880);
not NOT1 (N896, N894);
nand NAND4 (N897, N891, N652, N615, N402);
nor NOR4 (N898, N867, N502, N333, N451);
nand NAND4 (N899, N890, N53, N72, N825);
buf BUF1 (N900, N897);
nor NOR3 (N901, N899, N517, N46);
buf BUF1 (N902, N901);
nor NOR2 (N903, N902, N614);
nor NOR2 (N904, N900, N556);
nor NOR4 (N905, N903, N64, N801, N290);
buf BUF1 (N906, N893);
nand NAND3 (N907, N881, N223, N474);
buf BUF1 (N908, N896);
buf BUF1 (N909, N885);
buf BUF1 (N910, N905);
xor XOR2 (N911, N909, N157);
buf BUF1 (N912, N892);
or OR2 (N913, N912, N897);
not NOT1 (N914, N904);
xor XOR2 (N915, N911, N234);
buf BUF1 (N916, N907);
nand NAND2 (N917, N889, N204);
not NOT1 (N918, N906);
and AND3 (N919, N908, N259, N735);
or OR2 (N920, N910, N72);
and AND2 (N921, N915, N183);
nand NAND2 (N922, N898, N17);
nand NAND4 (N923, N919, N820, N744, N349);
nor NOR4 (N924, N895, N394, N97, N793);
or OR3 (N925, N916, N537, N479);
nand NAND3 (N926, N921, N874, N875);
or OR2 (N927, N923, N866);
buf BUF1 (N928, N917);
buf BUF1 (N929, N922);
and AND2 (N930, N928, N424);
and AND2 (N931, N918, N319);
not NOT1 (N932, N929);
and AND3 (N933, N914, N372, N266);
buf BUF1 (N934, N913);
and AND3 (N935, N931, N413, N670);
xor XOR2 (N936, N926, N928);
buf BUF1 (N937, N935);
nand NAND3 (N938, N932, N259, N116);
buf BUF1 (N939, N930);
not NOT1 (N940, N934);
buf BUF1 (N941, N925);
xor XOR2 (N942, N940, N885);
not NOT1 (N943, N941);
not NOT1 (N944, N943);
or OR4 (N945, N933, N574, N63, N223);
buf BUF1 (N946, N920);
nor NOR2 (N947, N939, N25);
nor NOR3 (N948, N936, N173, N349);
not NOT1 (N949, N937);
not NOT1 (N950, N949);
nor NOR2 (N951, N950, N918);
buf BUF1 (N952, N924);
xor XOR2 (N953, N938, N464);
not NOT1 (N954, N953);
and AND4 (N955, N951, N443, N192, N75);
xor XOR2 (N956, N948, N901);
not NOT1 (N957, N945);
not NOT1 (N958, N954);
or OR3 (N959, N946, N728, N806);
buf BUF1 (N960, N942);
xor XOR2 (N961, N947, N128);
not NOT1 (N962, N960);
xor XOR2 (N963, N959, N336);
buf BUF1 (N964, N957);
or OR2 (N965, N955, N700);
nor NOR2 (N966, N961, N319);
buf BUF1 (N967, N927);
not NOT1 (N968, N952);
xor XOR2 (N969, N956, N534);
nor NOR3 (N970, N964, N80, N132);
xor XOR2 (N971, N963, N608);
buf BUF1 (N972, N944);
buf BUF1 (N973, N971);
nand NAND2 (N974, N962, N84);
buf BUF1 (N975, N968);
and AND3 (N976, N973, N159, N175);
or OR4 (N977, N967, N480, N546, N49);
xor XOR2 (N978, N976, N183);
or OR2 (N979, N972, N829);
nand NAND4 (N980, N966, N331, N683, N817);
not NOT1 (N981, N975);
or OR4 (N982, N969, N522, N62, N557);
not NOT1 (N983, N974);
not NOT1 (N984, N977);
not NOT1 (N985, N983);
or OR2 (N986, N970, N749);
xor XOR2 (N987, N979, N433);
not NOT1 (N988, N965);
not NOT1 (N989, N980);
xor XOR2 (N990, N982, N896);
buf BUF1 (N991, N986);
nor NOR3 (N992, N958, N793, N990);
and AND3 (N993, N257, N340, N173);
buf BUF1 (N994, N988);
or OR4 (N995, N981, N881, N693, N246);
nand NAND3 (N996, N987, N763, N856);
and AND3 (N997, N992, N17, N927);
not NOT1 (N998, N993);
nor NOR4 (N999, N994, N656, N644, N257);
nor NOR4 (N1000, N984, N872, N837, N325);
xor XOR2 (N1001, N998, N491);
nand NAND3 (N1002, N1000, N748, N363);
not NOT1 (N1003, N989);
nand NAND2 (N1004, N991, N681);
buf BUF1 (N1005, N985);
or OR4 (N1006, N978, N509, N419, N382);
not NOT1 (N1007, N997);
and AND4 (N1008, N1006, N677, N603, N694);
or OR2 (N1009, N1001, N797);
nand NAND2 (N1010, N1004, N103);
buf BUF1 (N1011, N1010);
xor XOR2 (N1012, N1009, N513);
nand NAND2 (N1013, N996, N771);
nor NOR4 (N1014, N1013, N912, N355, N456);
or OR2 (N1015, N1002, N65);
and AND4 (N1016, N1014, N891, N569, N694);
and AND2 (N1017, N1012, N764);
nor NOR2 (N1018, N1005, N456);
or OR4 (N1019, N1017, N297, N188, N860);
xor XOR2 (N1020, N1011, N980);
buf BUF1 (N1021, N1015);
xor XOR2 (N1022, N1019, N706);
and AND4 (N1023, N1018, N612, N364, N674);
or OR4 (N1024, N999, N317, N243, N318);
not NOT1 (N1025, N1007);
buf BUF1 (N1026, N1003);
and AND2 (N1027, N1008, N475);
not NOT1 (N1028, N1027);
and AND4 (N1029, N1024, N293, N32, N445);
xor XOR2 (N1030, N1029, N603);
xor XOR2 (N1031, N995, N508);
nand NAND2 (N1032, N1028, N952);
nor NOR4 (N1033, N1031, N933, N933, N832);
or OR3 (N1034, N1033, N272, N527);
xor XOR2 (N1035, N1030, N825);
or OR3 (N1036, N1032, N709, N272);
buf BUF1 (N1037, N1016);
buf BUF1 (N1038, N1025);
nand NAND3 (N1039, N1035, N995, N416);
nand NAND2 (N1040, N1039, N256);
buf BUF1 (N1041, N1036);
nor NOR4 (N1042, N1041, N434, N601, N797);
xor XOR2 (N1043, N1020, N178);
buf BUF1 (N1044, N1040);
nand NAND2 (N1045, N1044, N735);
buf BUF1 (N1046, N1022);
and AND2 (N1047, N1034, N101);
nand NAND2 (N1048, N1047, N416);
nor NOR3 (N1049, N1043, N973, N601);
and AND4 (N1050, N1042, N454, N110, N43);
buf BUF1 (N1051, N1045);
xor XOR2 (N1052, N1050, N710);
nand NAND3 (N1053, N1021, N825, N673);
xor XOR2 (N1054, N1037, N691);
not NOT1 (N1055, N1049);
not NOT1 (N1056, N1053);
and AND2 (N1057, N1038, N707);
and AND2 (N1058, N1026, N400);
nor NOR4 (N1059, N1052, N835, N164, N338);
buf BUF1 (N1060, N1055);
buf BUF1 (N1061, N1057);
or OR2 (N1062, N1023, N861);
or OR3 (N1063, N1051, N96, N629);
nor NOR2 (N1064, N1059, N297);
nand NAND2 (N1065, N1046, N502);
or OR4 (N1066, N1063, N820, N430, N302);
not NOT1 (N1067, N1056);
buf BUF1 (N1068, N1054);
not NOT1 (N1069, N1067);
or OR2 (N1070, N1066, N251);
nand NAND4 (N1071, N1062, N933, N871, N8);
buf BUF1 (N1072, N1064);
buf BUF1 (N1073, N1071);
nor NOR4 (N1074, N1072, N265, N269, N19);
xor XOR2 (N1075, N1058, N965);
nor NOR2 (N1076, N1061, N361);
xor XOR2 (N1077, N1075, N932);
nand NAND3 (N1078, N1048, N607, N364);
nor NOR2 (N1079, N1074, N284);
buf BUF1 (N1080, N1073);
not NOT1 (N1081, N1078);
not NOT1 (N1082, N1080);
buf BUF1 (N1083, N1082);
buf BUF1 (N1084, N1081);
and AND3 (N1085, N1084, N743, N441);
nor NOR3 (N1086, N1069, N333, N210);
xor XOR2 (N1087, N1065, N647);
buf BUF1 (N1088, N1070);
xor XOR2 (N1089, N1087, N91);
or OR2 (N1090, N1085, N738);
or OR3 (N1091, N1077, N199, N580);
xor XOR2 (N1092, N1090, N975);
nor NOR4 (N1093, N1086, N693, N718, N160);
nor NOR3 (N1094, N1079, N300, N242);
buf BUF1 (N1095, N1094);
and AND3 (N1096, N1068, N728, N814);
or OR3 (N1097, N1083, N937, N831);
not NOT1 (N1098, N1095);
nand NAND3 (N1099, N1092, N402, N38);
buf BUF1 (N1100, N1076);
nand NAND4 (N1101, N1060, N451, N339, N302);
not NOT1 (N1102, N1088);
or OR4 (N1103, N1102, N1022, N705, N469);
not NOT1 (N1104, N1101);
and AND3 (N1105, N1103, N284, N657);
nor NOR3 (N1106, N1099, N604, N77);
nor NOR3 (N1107, N1100, N848, N554);
and AND3 (N1108, N1105, N751, N484);
nand NAND3 (N1109, N1108, N425, N119);
xor XOR2 (N1110, N1091, N943);
nand NAND3 (N1111, N1107, N493, N367);
buf BUF1 (N1112, N1089);
nor NOR3 (N1113, N1104, N584, N517);
buf BUF1 (N1114, N1093);
not NOT1 (N1115, N1098);
xor XOR2 (N1116, N1115, N17);
buf BUF1 (N1117, N1113);
or OR4 (N1118, N1111, N748, N230, N892);
buf BUF1 (N1119, N1110);
and AND2 (N1120, N1097, N414);
buf BUF1 (N1121, N1109);
xor XOR2 (N1122, N1096, N61);
nand NAND4 (N1123, N1112, N392, N1013, N518);
or OR2 (N1124, N1118, N828);
and AND2 (N1125, N1106, N767);
xor XOR2 (N1126, N1122, N920);
and AND3 (N1127, N1117, N524, N453);
nand NAND4 (N1128, N1120, N163, N605, N349);
nand NAND4 (N1129, N1128, N237, N877, N1054);
nand NAND2 (N1130, N1126, N335);
not NOT1 (N1131, N1123);
or OR3 (N1132, N1114, N981, N174);
and AND4 (N1133, N1125, N994, N748, N965);
nand NAND2 (N1134, N1121, N632);
or OR2 (N1135, N1133, N973);
buf BUF1 (N1136, N1130);
and AND2 (N1137, N1136, N1108);
nor NOR3 (N1138, N1127, N599, N664);
nand NAND2 (N1139, N1124, N664);
nor NOR3 (N1140, N1119, N704, N556);
nand NAND4 (N1141, N1135, N350, N719, N160);
buf BUF1 (N1142, N1138);
buf BUF1 (N1143, N1129);
not NOT1 (N1144, N1134);
nor NOR3 (N1145, N1137, N298, N503);
or OR4 (N1146, N1116, N915, N534, N328);
or OR4 (N1147, N1143, N51, N748, N639);
nand NAND4 (N1148, N1140, N773, N114, N657);
or OR3 (N1149, N1146, N284, N832);
nand NAND3 (N1150, N1147, N7, N430);
or OR3 (N1151, N1148, N93, N966);
nand NAND3 (N1152, N1145, N285, N966);
not NOT1 (N1153, N1142);
and AND4 (N1154, N1152, N227, N1152, N760);
not NOT1 (N1155, N1150);
and AND3 (N1156, N1132, N67, N379);
buf BUF1 (N1157, N1153);
nand NAND2 (N1158, N1131, N761);
or OR4 (N1159, N1144, N590, N396, N607);
xor XOR2 (N1160, N1139, N886);
buf BUF1 (N1161, N1155);
nor NOR4 (N1162, N1156, N1010, N813, N316);
not NOT1 (N1163, N1161);
xor XOR2 (N1164, N1162, N325);
nand NAND3 (N1165, N1141, N448, N154);
or OR2 (N1166, N1160, N828);
nor NOR2 (N1167, N1166, N771);
nand NAND3 (N1168, N1165, N101, N53);
not NOT1 (N1169, N1151);
or OR3 (N1170, N1167, N786, N1117);
nor NOR2 (N1171, N1159, N418);
xor XOR2 (N1172, N1168, N949);
xor XOR2 (N1173, N1157, N266);
buf BUF1 (N1174, N1149);
or OR3 (N1175, N1154, N409, N239);
or OR3 (N1176, N1173, N881, N231);
nor NOR2 (N1177, N1158, N773);
not NOT1 (N1178, N1175);
buf BUF1 (N1179, N1164);
nor NOR4 (N1180, N1172, N1127, N928, N479);
not NOT1 (N1181, N1177);
nand NAND2 (N1182, N1171, N449);
buf BUF1 (N1183, N1176);
buf BUF1 (N1184, N1163);
not NOT1 (N1185, N1181);
nand NAND2 (N1186, N1182, N722);
nand NAND2 (N1187, N1169, N64);
nand NAND2 (N1188, N1174, N750);
nand NAND4 (N1189, N1184, N450, N343, N1007);
buf BUF1 (N1190, N1170);
nor NOR2 (N1191, N1179, N573);
xor XOR2 (N1192, N1183, N264);
nand NAND2 (N1193, N1189, N599);
or OR2 (N1194, N1178, N395);
xor XOR2 (N1195, N1191, N967);
not NOT1 (N1196, N1187);
nor NOR2 (N1197, N1196, N353);
or OR3 (N1198, N1186, N627, N918);
or OR2 (N1199, N1188, N579);
buf BUF1 (N1200, N1199);
not NOT1 (N1201, N1193);
xor XOR2 (N1202, N1194, N552);
xor XOR2 (N1203, N1201, N111);
xor XOR2 (N1204, N1180, N723);
nand NAND4 (N1205, N1200, N673, N622, N646);
xor XOR2 (N1206, N1198, N221);
xor XOR2 (N1207, N1203, N719);
or OR3 (N1208, N1197, N193, N386);
or OR4 (N1209, N1204, N601, N812, N713);
not NOT1 (N1210, N1185);
nand NAND3 (N1211, N1202, N718, N307);
not NOT1 (N1212, N1205);
buf BUF1 (N1213, N1207);
nand NAND3 (N1214, N1213, N233, N1111);
not NOT1 (N1215, N1195);
or OR2 (N1216, N1192, N1028);
and AND4 (N1217, N1216, N946, N782, N216);
or OR4 (N1218, N1214, N238, N999, N283);
nor NOR4 (N1219, N1218, N338, N481, N424);
buf BUF1 (N1220, N1210);
nand NAND3 (N1221, N1212, N987, N952);
xor XOR2 (N1222, N1217, N618);
nor NOR3 (N1223, N1211, N236, N80);
or OR3 (N1224, N1208, N1065, N258);
nand NAND4 (N1225, N1222, N819, N289, N651);
buf BUF1 (N1226, N1219);
and AND4 (N1227, N1226, N685, N680, N444);
nand NAND3 (N1228, N1227, N376, N773);
nor NOR2 (N1229, N1225, N786);
nand NAND2 (N1230, N1221, N562);
not NOT1 (N1231, N1190);
nand NAND4 (N1232, N1231, N300, N390, N641);
not NOT1 (N1233, N1228);
and AND4 (N1234, N1232, N1010, N361, N404);
buf BUF1 (N1235, N1224);
nor NOR3 (N1236, N1209, N1191, N428);
or OR2 (N1237, N1223, N566);
not NOT1 (N1238, N1215);
xor XOR2 (N1239, N1220, N1087);
nand NAND2 (N1240, N1236, N957);
buf BUF1 (N1241, N1233);
nor NOR4 (N1242, N1230, N916, N670, N648);
nor NOR3 (N1243, N1234, N246, N619);
xor XOR2 (N1244, N1238, N733);
buf BUF1 (N1245, N1237);
nor NOR4 (N1246, N1229, N174, N707, N245);
nor NOR2 (N1247, N1206, N276);
buf BUF1 (N1248, N1246);
or OR3 (N1249, N1239, N959, N259);
and AND2 (N1250, N1247, N898);
buf BUF1 (N1251, N1245);
not NOT1 (N1252, N1248);
buf BUF1 (N1253, N1240);
buf BUF1 (N1254, N1242);
buf BUF1 (N1255, N1241);
not NOT1 (N1256, N1235);
and AND3 (N1257, N1249, N501, N791);
xor XOR2 (N1258, N1254, N583);
buf BUF1 (N1259, N1253);
not NOT1 (N1260, N1243);
and AND3 (N1261, N1250, N236, N802);
nand NAND2 (N1262, N1260, N639);
nand NAND4 (N1263, N1257, N609, N857, N515);
xor XOR2 (N1264, N1251, N178);
and AND3 (N1265, N1259, N897, N1020);
nand NAND4 (N1266, N1264, N1130, N96, N190);
not NOT1 (N1267, N1262);
and AND2 (N1268, N1267, N767);
and AND3 (N1269, N1256, N1142, N985);
and AND2 (N1270, N1252, N181);
or OR3 (N1271, N1265, N506, N556);
buf BUF1 (N1272, N1263);
nor NOR4 (N1273, N1268, N402, N959, N1253);
nand NAND3 (N1274, N1269, N374, N734);
nand NAND3 (N1275, N1273, N1114, N194);
buf BUF1 (N1276, N1244);
nor NOR3 (N1277, N1270, N219, N289);
xor XOR2 (N1278, N1275, N568);
or OR4 (N1279, N1274, N592, N960, N188);
not NOT1 (N1280, N1261);
and AND2 (N1281, N1258, N1075);
buf BUF1 (N1282, N1276);
xor XOR2 (N1283, N1280, N404);
xor XOR2 (N1284, N1282, N926);
nor NOR3 (N1285, N1277, N248, N612);
or OR3 (N1286, N1271, N348, N95);
or OR3 (N1287, N1278, N598, N361);
not NOT1 (N1288, N1279);
buf BUF1 (N1289, N1287);
and AND2 (N1290, N1284, N1158);
and AND4 (N1291, N1290, N787, N467, N664);
xor XOR2 (N1292, N1291, N24);
buf BUF1 (N1293, N1286);
and AND2 (N1294, N1272, N931);
nor NOR4 (N1295, N1285, N672, N226, N365);
and AND4 (N1296, N1283, N1222, N939, N572);
and AND2 (N1297, N1281, N976);
nor NOR2 (N1298, N1295, N774);
buf BUF1 (N1299, N1294);
xor XOR2 (N1300, N1293, N1023);
buf BUF1 (N1301, N1266);
buf BUF1 (N1302, N1296);
not NOT1 (N1303, N1289);
or OR4 (N1304, N1300, N626, N571, N600);
or OR2 (N1305, N1302, N1001);
nand NAND4 (N1306, N1292, N168, N423, N274);
not NOT1 (N1307, N1255);
nor NOR4 (N1308, N1301, N288, N263, N223);
nor NOR3 (N1309, N1298, N920, N64);
nand NAND2 (N1310, N1303, N806);
buf BUF1 (N1311, N1288);
xor XOR2 (N1312, N1310, N1164);
and AND4 (N1313, N1306, N454, N571, N464);
nand NAND4 (N1314, N1313, N1226, N597, N1213);
xor XOR2 (N1315, N1312, N685);
nor NOR3 (N1316, N1308, N779, N473);
and AND4 (N1317, N1307, N1192, N821, N235);
xor XOR2 (N1318, N1305, N779);
xor XOR2 (N1319, N1318, N919);
xor XOR2 (N1320, N1299, N1319);
and AND4 (N1321, N421, N703, N1227, N1070);
or OR2 (N1322, N1304, N997);
and AND2 (N1323, N1311, N21);
buf BUF1 (N1324, N1314);
xor XOR2 (N1325, N1324, N543);
buf BUF1 (N1326, N1309);
nand NAND3 (N1327, N1320, N454, N17);
buf BUF1 (N1328, N1326);
xor XOR2 (N1329, N1325, N293);
buf BUF1 (N1330, N1327);
nand NAND2 (N1331, N1317, N1245);
and AND4 (N1332, N1297, N561, N365, N491);
nor NOR2 (N1333, N1328, N134);
nand NAND2 (N1334, N1323, N217);
nor NOR3 (N1335, N1322, N358, N835);
xor XOR2 (N1336, N1321, N1230);
nand NAND4 (N1337, N1334, N884, N112, N196);
or OR3 (N1338, N1333, N1219, N1055);
and AND2 (N1339, N1331, N1057);
xor XOR2 (N1340, N1332, N1050);
and AND3 (N1341, N1335, N4, N1259);
nor NOR2 (N1342, N1330, N191);
buf BUF1 (N1343, N1341);
nand NAND3 (N1344, N1340, N1185, N205);
nand NAND2 (N1345, N1329, N894);
and AND2 (N1346, N1345, N969);
xor XOR2 (N1347, N1315, N565);
nor NOR2 (N1348, N1342, N1219);
and AND2 (N1349, N1339, N1178);
xor XOR2 (N1350, N1344, N586);
or OR2 (N1351, N1337, N37);
nand NAND4 (N1352, N1316, N676, N110, N944);
buf BUF1 (N1353, N1347);
and AND3 (N1354, N1346, N272, N1012);
not NOT1 (N1355, N1354);
or OR3 (N1356, N1351, N382, N952);
not NOT1 (N1357, N1348);
buf BUF1 (N1358, N1357);
buf BUF1 (N1359, N1353);
or OR3 (N1360, N1338, N1165, N411);
nand NAND2 (N1361, N1356, N1012);
xor XOR2 (N1362, N1355, N259);
nor NOR3 (N1363, N1361, N366, N636);
buf BUF1 (N1364, N1363);
buf BUF1 (N1365, N1349);
and AND2 (N1366, N1350, N67);
not NOT1 (N1367, N1362);
buf BUF1 (N1368, N1343);
xor XOR2 (N1369, N1360, N1217);
nor NOR4 (N1370, N1358, N1308, N1333, N18);
xor XOR2 (N1371, N1368, N1307);
buf BUF1 (N1372, N1359);
nand NAND3 (N1373, N1369, N1326, N1064);
buf BUF1 (N1374, N1371);
buf BUF1 (N1375, N1365);
not NOT1 (N1376, N1372);
buf BUF1 (N1377, N1364);
or OR2 (N1378, N1374, N102);
nand NAND3 (N1379, N1367, N1201, N119);
not NOT1 (N1380, N1377);
not NOT1 (N1381, N1336);
and AND4 (N1382, N1370, N1243, N841, N230);
nor NOR4 (N1383, N1382, N437, N941, N1068);
xor XOR2 (N1384, N1381, N30);
buf BUF1 (N1385, N1379);
not NOT1 (N1386, N1383);
nor NOR2 (N1387, N1373, N1176);
xor XOR2 (N1388, N1378, N240);
and AND3 (N1389, N1384, N860, N383);
nand NAND4 (N1390, N1352, N1343, N100, N810);
nor NOR3 (N1391, N1388, N962, N248);
nand NAND2 (N1392, N1385, N1281);
nor NOR3 (N1393, N1392, N154, N429);
nand NAND3 (N1394, N1366, N847, N985);
xor XOR2 (N1395, N1387, N1161);
xor XOR2 (N1396, N1386, N1358);
nand NAND3 (N1397, N1390, N668, N1230);
nor NOR2 (N1398, N1389, N1177);
xor XOR2 (N1399, N1393, N330);
xor XOR2 (N1400, N1399, N1158);
buf BUF1 (N1401, N1376);
xor XOR2 (N1402, N1396, N543);
and AND2 (N1403, N1400, N901);
or OR4 (N1404, N1402, N849, N1040, N118);
nor NOR2 (N1405, N1401, N509);
nor NOR3 (N1406, N1397, N198, N976);
and AND2 (N1407, N1391, N103);
nand NAND2 (N1408, N1406, N286);
xor XOR2 (N1409, N1375, N941);
nor NOR4 (N1410, N1407, N25, N725, N1095);
and AND4 (N1411, N1404, N246, N1342, N863);
or OR2 (N1412, N1398, N701);
buf BUF1 (N1413, N1410);
buf BUF1 (N1414, N1412);
nor NOR2 (N1415, N1413, N1123);
xor XOR2 (N1416, N1395, N1160);
nand NAND4 (N1417, N1408, N1355, N33, N470);
or OR2 (N1418, N1417, N17);
xor XOR2 (N1419, N1418, N374);
nor NOR2 (N1420, N1419, N424);
not NOT1 (N1421, N1416);
buf BUF1 (N1422, N1403);
not NOT1 (N1423, N1411);
not NOT1 (N1424, N1414);
or OR3 (N1425, N1422, N1189, N777);
nor NOR2 (N1426, N1425, N393);
buf BUF1 (N1427, N1423);
not NOT1 (N1428, N1420);
not NOT1 (N1429, N1424);
not NOT1 (N1430, N1421);
or OR3 (N1431, N1380, N930, N364);
nand NAND3 (N1432, N1431, N733, N553);
not NOT1 (N1433, N1394);
or OR3 (N1434, N1433, N911, N1084);
xor XOR2 (N1435, N1409, N493);
not NOT1 (N1436, N1428);
nor NOR2 (N1437, N1415, N1319);
nand NAND2 (N1438, N1427, N148);
nand NAND3 (N1439, N1435, N625, N1133);
or OR2 (N1440, N1429, N16);
and AND2 (N1441, N1432, N1080);
nor NOR2 (N1442, N1441, N1376);
nor NOR4 (N1443, N1430, N781, N1426, N1438);
nor NOR3 (N1444, N46, N293, N354);
nand NAND3 (N1445, N1167, N1016, N1036);
not NOT1 (N1446, N1434);
nand NAND4 (N1447, N1446, N1169, N1306, N1238);
or OR3 (N1448, N1440, N29, N1006);
and AND4 (N1449, N1437, N980, N933, N340);
nor NOR2 (N1450, N1436, N627);
and AND2 (N1451, N1439, N423);
buf BUF1 (N1452, N1444);
nand NAND3 (N1453, N1447, N1309, N1231);
xor XOR2 (N1454, N1448, N832);
nor NOR4 (N1455, N1451, N463, N108, N260);
buf BUF1 (N1456, N1405);
nand NAND3 (N1457, N1449, N437, N1229);
nor NOR4 (N1458, N1450, N1117, N1034, N1171);
or OR4 (N1459, N1457, N224, N198, N914);
xor XOR2 (N1460, N1458, N297);
xor XOR2 (N1461, N1454, N585);
and AND2 (N1462, N1453, N156);
not NOT1 (N1463, N1445);
buf BUF1 (N1464, N1442);
not NOT1 (N1465, N1443);
nand NAND4 (N1466, N1463, N983, N933, N946);
or OR3 (N1467, N1461, N12, N861);
nand NAND2 (N1468, N1467, N371);
buf BUF1 (N1469, N1459);
or OR2 (N1470, N1469, N1040);
and AND4 (N1471, N1456, N416, N1151, N655);
and AND4 (N1472, N1465, N73, N519, N828);
xor XOR2 (N1473, N1460, N1388);
or OR4 (N1474, N1468, N1396, N521, N526);
not NOT1 (N1475, N1455);
nor NOR4 (N1476, N1470, N500, N1443, N1251);
or OR4 (N1477, N1476, N1312, N587, N1362);
or OR4 (N1478, N1473, N743, N746, N1168);
xor XOR2 (N1479, N1462, N1419);
buf BUF1 (N1480, N1452);
xor XOR2 (N1481, N1475, N374);
nand NAND4 (N1482, N1466, N515, N113, N861);
nor NOR3 (N1483, N1471, N1181, N641);
not NOT1 (N1484, N1482);
and AND4 (N1485, N1464, N979, N499, N803);
buf BUF1 (N1486, N1474);
buf BUF1 (N1487, N1484);
or OR4 (N1488, N1478, N553, N344, N884);
nor NOR2 (N1489, N1479, N145);
and AND3 (N1490, N1483, N1043, N1359);
xor XOR2 (N1491, N1480, N188);
xor XOR2 (N1492, N1488, N273);
not NOT1 (N1493, N1492);
nand NAND4 (N1494, N1490, N684, N1338, N990);
nand NAND3 (N1495, N1491, N1394, N794);
and AND2 (N1496, N1495, N1451);
xor XOR2 (N1497, N1486, N627);
buf BUF1 (N1498, N1493);
buf BUF1 (N1499, N1498);
not NOT1 (N1500, N1487);
not NOT1 (N1501, N1500);
xor XOR2 (N1502, N1472, N1156);
not NOT1 (N1503, N1485);
or OR4 (N1504, N1494, N1047, N628, N577);
nor NOR3 (N1505, N1477, N451, N700);
nor NOR3 (N1506, N1502, N432, N1441);
or OR4 (N1507, N1489, N475, N120, N1112);
not NOT1 (N1508, N1501);
xor XOR2 (N1509, N1506, N423);
xor XOR2 (N1510, N1508, N32);
not NOT1 (N1511, N1505);
nor NOR4 (N1512, N1511, N681, N1050, N707);
nor NOR3 (N1513, N1499, N1264, N424);
buf BUF1 (N1514, N1507);
xor XOR2 (N1515, N1512, N974);
and AND4 (N1516, N1510, N468, N527, N1286);
nor NOR4 (N1517, N1504, N82, N266, N1359);
nor NOR4 (N1518, N1514, N743, N984, N1324);
not NOT1 (N1519, N1509);
nand NAND2 (N1520, N1518, N1037);
and AND4 (N1521, N1497, N1356, N590, N1499);
buf BUF1 (N1522, N1520);
nor NOR3 (N1523, N1496, N499, N727);
or OR3 (N1524, N1519, N728, N965);
and AND2 (N1525, N1481, N1168);
xor XOR2 (N1526, N1521, N771);
nor NOR4 (N1527, N1522, N525, N365, N1388);
and AND2 (N1528, N1517, N1264);
or OR3 (N1529, N1516, N948, N556);
buf BUF1 (N1530, N1513);
nand NAND2 (N1531, N1523, N305);
and AND2 (N1532, N1524, N247);
buf BUF1 (N1533, N1532);
xor XOR2 (N1534, N1530, N820);
nand NAND2 (N1535, N1534, N513);
or OR2 (N1536, N1503, N314);
xor XOR2 (N1537, N1528, N964);
or OR4 (N1538, N1527, N705, N729, N1323);
xor XOR2 (N1539, N1537, N1047);
and AND4 (N1540, N1536, N1424, N1047, N1093);
or OR4 (N1541, N1529, N1200, N898, N170);
buf BUF1 (N1542, N1525);
buf BUF1 (N1543, N1540);
or OR4 (N1544, N1538, N1366, N155, N1186);
buf BUF1 (N1545, N1539);
not NOT1 (N1546, N1542);
not NOT1 (N1547, N1535);
and AND3 (N1548, N1543, N714, N330);
or OR3 (N1549, N1533, N849, N1273);
nor NOR2 (N1550, N1526, N1197);
and AND2 (N1551, N1546, N1482);
and AND4 (N1552, N1531, N710, N251, N1294);
xor XOR2 (N1553, N1545, N260);
not NOT1 (N1554, N1552);
and AND2 (N1555, N1541, N871);
not NOT1 (N1556, N1554);
nand NAND3 (N1557, N1551, N543, N283);
or OR2 (N1558, N1515, N913);
nand NAND4 (N1559, N1544, N1115, N233, N792);
nor NOR2 (N1560, N1550, N1556);
not NOT1 (N1561, N1066);
nand NAND3 (N1562, N1547, N580, N1506);
or OR2 (N1563, N1555, N1440);
nand NAND4 (N1564, N1558, N960, N919, N1450);
or OR4 (N1565, N1563, N30, N1029, N562);
or OR3 (N1566, N1549, N330, N1142);
xor XOR2 (N1567, N1557, N858);
and AND4 (N1568, N1562, N509, N1297, N448);
and AND2 (N1569, N1566, N370);
buf BUF1 (N1570, N1548);
or OR2 (N1571, N1553, N1042);
buf BUF1 (N1572, N1567);
nand NAND4 (N1573, N1560, N891, N1515, N1476);
nor NOR2 (N1574, N1565, N542);
and AND4 (N1575, N1561, N84, N864, N212);
buf BUF1 (N1576, N1570);
nor NOR2 (N1577, N1559, N651);
not NOT1 (N1578, N1575);
nand NAND4 (N1579, N1576, N606, N1461, N634);
or OR3 (N1580, N1571, N1503, N1191);
not NOT1 (N1581, N1573);
xor XOR2 (N1582, N1569, N686);
nand NAND3 (N1583, N1581, N764, N25);
not NOT1 (N1584, N1568);
nand NAND4 (N1585, N1579, N80, N1568, N110);
nand NAND3 (N1586, N1564, N1347, N482);
nor NOR3 (N1587, N1586, N714, N1459);
nand NAND4 (N1588, N1582, N1073, N594, N1024);
or OR3 (N1589, N1578, N1093, N1342);
nand NAND4 (N1590, N1585, N475, N948, N854);
nor NOR3 (N1591, N1584, N115, N228);
nand NAND3 (N1592, N1588, N407, N311);
or OR2 (N1593, N1583, N1036);
buf BUF1 (N1594, N1591);
nor NOR3 (N1595, N1594, N150, N61);
nand NAND4 (N1596, N1593, N689, N446, N768);
buf BUF1 (N1597, N1574);
xor XOR2 (N1598, N1580, N987);
nand NAND3 (N1599, N1572, N1083, N309);
or OR4 (N1600, N1590, N643, N1157, N1426);
buf BUF1 (N1601, N1577);
or OR4 (N1602, N1589, N946, N922, N600);
or OR4 (N1603, N1599, N238, N788, N836);
buf BUF1 (N1604, N1597);
and AND2 (N1605, N1592, N509);
and AND2 (N1606, N1601, N1435);
or OR3 (N1607, N1605, N940, N961);
nor NOR2 (N1608, N1604, N1480);
not NOT1 (N1609, N1606);
and AND3 (N1610, N1602, N1526, N87);
and AND2 (N1611, N1600, N722);
xor XOR2 (N1612, N1608, N647);
not NOT1 (N1613, N1609);
buf BUF1 (N1614, N1612);
or OR4 (N1615, N1613, N643, N1052, N1195);
buf BUF1 (N1616, N1607);
not NOT1 (N1617, N1615);
nand NAND2 (N1618, N1614, N1568);
nor NOR2 (N1619, N1611, N1476);
nand NAND2 (N1620, N1618, N451);
buf BUF1 (N1621, N1619);
xor XOR2 (N1622, N1598, N1524);
and AND4 (N1623, N1616, N1182, N749, N618);
buf BUF1 (N1624, N1617);
and AND4 (N1625, N1623, N267, N647, N265);
nor NOR2 (N1626, N1610, N1359);
buf BUF1 (N1627, N1620);
and AND4 (N1628, N1622, N657, N1160, N61);
and AND3 (N1629, N1621, N948, N1357);
xor XOR2 (N1630, N1587, N713);
nor NOR3 (N1631, N1630, N13, N1337);
nand NAND2 (N1632, N1627, N569);
not NOT1 (N1633, N1628);
nor NOR4 (N1634, N1626, N755, N1020, N1047);
nand NAND4 (N1635, N1603, N1544, N136, N291);
not NOT1 (N1636, N1633);
and AND3 (N1637, N1595, N56, N680);
and AND3 (N1638, N1631, N1494, N1433);
xor XOR2 (N1639, N1634, N1506);
nor NOR2 (N1640, N1639, N198);
buf BUF1 (N1641, N1640);
and AND4 (N1642, N1636, N1332, N1591, N910);
nor NOR4 (N1643, N1624, N561, N229, N2);
or OR2 (N1644, N1638, N201);
not NOT1 (N1645, N1625);
nor NOR3 (N1646, N1637, N1412, N71);
and AND3 (N1647, N1642, N1359, N1546);
not NOT1 (N1648, N1645);
not NOT1 (N1649, N1644);
not NOT1 (N1650, N1635);
nor NOR2 (N1651, N1632, N939);
buf BUF1 (N1652, N1643);
nor NOR2 (N1653, N1651, N751);
nor NOR3 (N1654, N1647, N234, N604);
xor XOR2 (N1655, N1629, N491);
buf BUF1 (N1656, N1648);
xor XOR2 (N1657, N1654, N889);
or OR3 (N1658, N1653, N607, N866);
not NOT1 (N1659, N1652);
or OR3 (N1660, N1657, N349, N1214);
or OR3 (N1661, N1660, N343, N1413);
nor NOR2 (N1662, N1650, N1259);
xor XOR2 (N1663, N1646, N795);
not NOT1 (N1664, N1641);
buf BUF1 (N1665, N1664);
nor NOR4 (N1666, N1649, N1200, N1013, N1131);
not NOT1 (N1667, N1655);
and AND2 (N1668, N1663, N134);
buf BUF1 (N1669, N1668);
nand NAND3 (N1670, N1666, N437, N1190);
buf BUF1 (N1671, N1669);
nand NAND4 (N1672, N1661, N262, N862, N1161);
xor XOR2 (N1673, N1656, N1505);
not NOT1 (N1674, N1596);
buf BUF1 (N1675, N1662);
buf BUF1 (N1676, N1672);
or OR3 (N1677, N1674, N9, N335);
buf BUF1 (N1678, N1670);
xor XOR2 (N1679, N1659, N221);
not NOT1 (N1680, N1676);
nand NAND2 (N1681, N1665, N135);
not NOT1 (N1682, N1671);
nand NAND4 (N1683, N1680, N1198, N162, N347);
or OR2 (N1684, N1667, N1531);
nor NOR3 (N1685, N1675, N953, N237);
nor NOR2 (N1686, N1658, N324);
buf BUF1 (N1687, N1684);
xor XOR2 (N1688, N1673, N1055);
not NOT1 (N1689, N1678);
or OR2 (N1690, N1682, N263);
xor XOR2 (N1691, N1685, N1360);
and AND4 (N1692, N1688, N166, N1271, N1182);
buf BUF1 (N1693, N1681);
or OR2 (N1694, N1677, N222);
buf BUF1 (N1695, N1691);
nor NOR4 (N1696, N1690, N194, N1098, N1538);
xor XOR2 (N1697, N1693, N858);
buf BUF1 (N1698, N1689);
and AND4 (N1699, N1698, N849, N207, N230);
nand NAND4 (N1700, N1696, N326, N1421, N556);
not NOT1 (N1701, N1686);
buf BUF1 (N1702, N1695);
buf BUF1 (N1703, N1697);
or OR3 (N1704, N1692, N1171, N463);
and AND4 (N1705, N1700, N750, N597, N1273);
nand NAND4 (N1706, N1701, N1445, N477, N99);
xor XOR2 (N1707, N1703, N949);
nand NAND3 (N1708, N1704, N979, N1362);
nand NAND3 (N1709, N1708, N354, N355);
nand NAND4 (N1710, N1707, N1528, N1380, N84);
nand NAND4 (N1711, N1687, N1273, N747, N30);
nor NOR2 (N1712, N1699, N93);
nor NOR2 (N1713, N1706, N237);
nand NAND4 (N1714, N1710, N956, N705, N104);
and AND2 (N1715, N1683, N1528);
or OR2 (N1716, N1712, N741);
xor XOR2 (N1717, N1714, N58);
or OR3 (N1718, N1709, N120, N1212);
not NOT1 (N1719, N1713);
not NOT1 (N1720, N1702);
and AND3 (N1721, N1711, N220, N307);
buf BUF1 (N1722, N1716);
nand NAND2 (N1723, N1679, N1378);
xor XOR2 (N1724, N1715, N1212);
xor XOR2 (N1725, N1722, N176);
and AND3 (N1726, N1719, N610, N411);
xor XOR2 (N1727, N1725, N827);
not NOT1 (N1728, N1694);
nor NOR2 (N1729, N1727, N930);
xor XOR2 (N1730, N1729, N97);
or OR2 (N1731, N1721, N3);
nand NAND2 (N1732, N1726, N1552);
buf BUF1 (N1733, N1728);
nand NAND4 (N1734, N1705, N954, N924, N675);
buf BUF1 (N1735, N1730);
nand NAND4 (N1736, N1723, N588, N752, N1120);
not NOT1 (N1737, N1736);
nand NAND2 (N1738, N1718, N442);
xor XOR2 (N1739, N1732, N818);
nor NOR4 (N1740, N1724, N874, N994, N1533);
nor NOR3 (N1741, N1731, N783, N351);
xor XOR2 (N1742, N1735, N543);
and AND3 (N1743, N1717, N1159, N1323);
or OR2 (N1744, N1740, N1519);
and AND2 (N1745, N1739, N852);
not NOT1 (N1746, N1743);
buf BUF1 (N1747, N1746);
or OR2 (N1748, N1720, N1523);
xor XOR2 (N1749, N1733, N1729);
nor NOR4 (N1750, N1749, N776, N238, N1300);
or OR2 (N1751, N1741, N1529);
nand NAND4 (N1752, N1750, N1004, N1627, N1656);
buf BUF1 (N1753, N1742);
or OR2 (N1754, N1751, N336);
xor XOR2 (N1755, N1754, N1467);
nand NAND2 (N1756, N1745, N45);
not NOT1 (N1757, N1747);
nand NAND3 (N1758, N1748, N803, N319);
nand NAND3 (N1759, N1753, N191, N981);
nor NOR3 (N1760, N1755, N137, N1038);
or OR3 (N1761, N1759, N851, N1566);
or OR3 (N1762, N1761, N1601, N370);
buf BUF1 (N1763, N1734);
not NOT1 (N1764, N1756);
and AND2 (N1765, N1744, N1121);
and AND2 (N1766, N1765, N1110);
nand NAND3 (N1767, N1738, N199, N706);
and AND3 (N1768, N1763, N1265, N1588);
nand NAND2 (N1769, N1757, N507);
nand NAND3 (N1770, N1760, N656, N572);
xor XOR2 (N1771, N1764, N852);
not NOT1 (N1772, N1769);
nand NAND2 (N1773, N1771, N1266);
or OR3 (N1774, N1768, N523, N801);
not NOT1 (N1775, N1773);
buf BUF1 (N1776, N1758);
and AND2 (N1777, N1737, N1557);
and AND4 (N1778, N1772, N800, N364, N1504);
xor XOR2 (N1779, N1777, N1286);
buf BUF1 (N1780, N1776);
or OR3 (N1781, N1762, N1724, N1403);
not NOT1 (N1782, N1766);
or OR3 (N1783, N1767, N925, N248);
nor NOR4 (N1784, N1752, N1734, N1296, N1135);
nor NOR3 (N1785, N1784, N921, N22);
not NOT1 (N1786, N1783);
and AND3 (N1787, N1774, N13, N299);
not NOT1 (N1788, N1782);
xor XOR2 (N1789, N1786, N1154);
nand NAND2 (N1790, N1770, N696);
or OR4 (N1791, N1785, N580, N1239, N226);
nand NAND3 (N1792, N1779, N311, N116);
xor XOR2 (N1793, N1775, N1239);
xor XOR2 (N1794, N1791, N1486);
or OR3 (N1795, N1793, N449, N631);
or OR2 (N1796, N1778, N1299);
not NOT1 (N1797, N1796);
nor NOR4 (N1798, N1788, N800, N1574, N441);
nand NAND4 (N1799, N1794, N404, N607, N1751);
and AND2 (N1800, N1787, N1324);
xor XOR2 (N1801, N1795, N1671);
not NOT1 (N1802, N1797);
buf BUF1 (N1803, N1801);
nor NOR2 (N1804, N1790, N106);
nand NAND3 (N1805, N1800, N1743, N884);
not NOT1 (N1806, N1792);
buf BUF1 (N1807, N1802);
xor XOR2 (N1808, N1804, N320);
and AND3 (N1809, N1805, N547, N1049);
nor NOR4 (N1810, N1803, N1809, N635, N810);
nor NOR4 (N1811, N643, N657, N1666, N800);
not NOT1 (N1812, N1806);
xor XOR2 (N1813, N1808, N1530);
xor XOR2 (N1814, N1780, N1129);
nand NAND2 (N1815, N1798, N1571);
not NOT1 (N1816, N1789);
buf BUF1 (N1817, N1814);
buf BUF1 (N1818, N1811);
xor XOR2 (N1819, N1818, N989);
xor XOR2 (N1820, N1813, N278);
xor XOR2 (N1821, N1807, N1819);
buf BUF1 (N1822, N1373);
nor NOR4 (N1823, N1817, N1131, N1612, N1591);
and AND3 (N1824, N1810, N1096, N1514);
or OR3 (N1825, N1821, N66, N330);
not NOT1 (N1826, N1816);
xor XOR2 (N1827, N1826, N1062);
not NOT1 (N1828, N1827);
xor XOR2 (N1829, N1781, N255);
or OR4 (N1830, N1829, N457, N141, N1806);
and AND4 (N1831, N1812, N840, N330, N330);
or OR2 (N1832, N1822, N1041);
not NOT1 (N1833, N1828);
and AND3 (N1834, N1820, N440, N29);
or OR4 (N1835, N1799, N37, N633, N1785);
buf BUF1 (N1836, N1832);
xor XOR2 (N1837, N1815, N1719);
buf BUF1 (N1838, N1835);
or OR4 (N1839, N1823, N675, N1516, N1384);
nand NAND4 (N1840, N1837, N1274, N426, N964);
and AND3 (N1841, N1834, N1234, N744);
xor XOR2 (N1842, N1840, N891);
xor XOR2 (N1843, N1838, N949);
nand NAND2 (N1844, N1836, N237);
buf BUF1 (N1845, N1842);
xor XOR2 (N1846, N1831, N306);
and AND4 (N1847, N1841, N632, N3, N1287);
nor NOR4 (N1848, N1839, N1090, N792, N1013);
xor XOR2 (N1849, N1846, N785);
nor NOR4 (N1850, N1825, N940, N1230, N1080);
xor XOR2 (N1851, N1830, N1034);
nor NOR3 (N1852, N1845, N672, N1337);
nand NAND3 (N1853, N1847, N730, N1266);
nor NOR2 (N1854, N1848, N1004);
nand NAND3 (N1855, N1850, N529, N401);
nor NOR4 (N1856, N1851, N1495, N1188, N1222);
or OR4 (N1857, N1855, N790, N217, N466);
xor XOR2 (N1858, N1824, N1561);
buf BUF1 (N1859, N1854);
buf BUF1 (N1860, N1843);
nor NOR2 (N1861, N1859, N92);
or OR4 (N1862, N1852, N1520, N939, N49);
buf BUF1 (N1863, N1849);
nor NOR3 (N1864, N1863, N1829, N632);
buf BUF1 (N1865, N1862);
nor NOR3 (N1866, N1861, N360, N687);
or OR2 (N1867, N1857, N903);
buf BUF1 (N1868, N1833);
or OR3 (N1869, N1865, N1643, N1575);
and AND3 (N1870, N1853, N1473, N1562);
or OR3 (N1871, N1860, N779, N1799);
or OR2 (N1872, N1844, N1408);
not NOT1 (N1873, N1856);
not NOT1 (N1874, N1868);
buf BUF1 (N1875, N1874);
and AND2 (N1876, N1871, N1653);
or OR4 (N1877, N1864, N553, N335, N1817);
nor NOR3 (N1878, N1870, N541, N1768);
buf BUF1 (N1879, N1858);
not NOT1 (N1880, N1875);
not NOT1 (N1881, N1876);
not NOT1 (N1882, N1878);
nand NAND3 (N1883, N1873, N1271, N28);
and AND4 (N1884, N1877, N734, N66, N1596);
nor NOR2 (N1885, N1866, N27);
nor NOR3 (N1886, N1884, N1652, N763);
or OR2 (N1887, N1881, N1614);
and AND2 (N1888, N1883, N795);
nor NOR4 (N1889, N1888, N989, N1869, N476);
nand NAND3 (N1890, N795, N550, N1345);
and AND3 (N1891, N1885, N1315, N17);
buf BUF1 (N1892, N1890);
not NOT1 (N1893, N1882);
xor XOR2 (N1894, N1892, N772);
or OR3 (N1895, N1889, N598, N1259);
or OR4 (N1896, N1893, N1888, N1564, N128);
buf BUF1 (N1897, N1895);
nand NAND3 (N1898, N1896, N1022, N441);
not NOT1 (N1899, N1886);
nor NOR3 (N1900, N1880, N1808, N1898);
buf BUF1 (N1901, N403);
xor XOR2 (N1902, N1894, N273);
buf BUF1 (N1903, N1867);
nor NOR3 (N1904, N1902, N114, N668);
buf BUF1 (N1905, N1879);
nor NOR3 (N1906, N1904, N649, N745);
not NOT1 (N1907, N1905);
xor XOR2 (N1908, N1897, N163);
and AND2 (N1909, N1872, N1101);
xor XOR2 (N1910, N1908, N1410);
xor XOR2 (N1911, N1909, N1432);
xor XOR2 (N1912, N1910, N100);
buf BUF1 (N1913, N1906);
or OR4 (N1914, N1913, N1584, N1534, N691);
nand NAND3 (N1915, N1911, N1558, N867);
nand NAND4 (N1916, N1912, N704, N1173, N1813);
buf BUF1 (N1917, N1907);
or OR2 (N1918, N1915, N1440);
and AND3 (N1919, N1918, N320, N372);
buf BUF1 (N1920, N1916);
or OR4 (N1921, N1903, N875, N1607, N206);
buf BUF1 (N1922, N1891);
nor NOR4 (N1923, N1922, N1190, N797, N694);
or OR3 (N1924, N1923, N1730, N1805);
and AND3 (N1925, N1887, N1276, N1356);
not NOT1 (N1926, N1914);
nand NAND3 (N1927, N1926, N680, N331);
and AND2 (N1928, N1900, N937);
and AND3 (N1929, N1917, N167, N1501);
and AND2 (N1930, N1924, N105);
xor XOR2 (N1931, N1929, N730);
nor NOR3 (N1932, N1930, N341, N1720);
or OR4 (N1933, N1931, N626, N1330, N268);
and AND2 (N1934, N1925, N1413);
nor NOR3 (N1935, N1927, N800, N673);
buf BUF1 (N1936, N1899);
or OR4 (N1937, N1919, N489, N521, N1016);
or OR2 (N1938, N1932, N30);
nor NOR3 (N1939, N1937, N1498, N435);
nor NOR3 (N1940, N1936, N1169, N885);
and AND3 (N1941, N1934, N567, N412);
not NOT1 (N1942, N1940);
nand NAND2 (N1943, N1941, N572);
xor XOR2 (N1944, N1920, N1078);
and AND4 (N1945, N1921, N1098, N1771, N16);
not NOT1 (N1946, N1942);
xor XOR2 (N1947, N1901, N1399);
buf BUF1 (N1948, N1944);
and AND2 (N1949, N1943, N162);
xor XOR2 (N1950, N1938, N1559);
xor XOR2 (N1951, N1948, N1574);
nand NAND3 (N1952, N1949, N1751, N573);
not NOT1 (N1953, N1928);
not NOT1 (N1954, N1953);
nand NAND4 (N1955, N1952, N418, N977, N1086);
and AND3 (N1956, N1933, N1312, N1164);
not NOT1 (N1957, N1947);
and AND3 (N1958, N1945, N292, N575);
not NOT1 (N1959, N1946);
xor XOR2 (N1960, N1954, N1435);
not NOT1 (N1961, N1959);
not NOT1 (N1962, N1957);
xor XOR2 (N1963, N1955, N188);
not NOT1 (N1964, N1960);
buf BUF1 (N1965, N1961);
nand NAND3 (N1966, N1962, N1345, N1646);
nor NOR4 (N1967, N1958, N1739, N549, N875);
xor XOR2 (N1968, N1939, N544);
nand NAND3 (N1969, N1956, N28, N1804);
buf BUF1 (N1970, N1935);
or OR3 (N1971, N1967, N1220, N1758);
not NOT1 (N1972, N1969);
not NOT1 (N1973, N1964);
nor NOR4 (N1974, N1963, N329, N1099, N1756);
nand NAND3 (N1975, N1950, N1598, N1324);
nand NAND2 (N1976, N1975, N483);
nor NOR3 (N1977, N1966, N311, N1555);
or OR4 (N1978, N1970, N1797, N1319, N1197);
and AND4 (N1979, N1972, N443, N880, N1804);
nand NAND4 (N1980, N1971, N341, N1758, N376);
and AND4 (N1981, N1974, N1062, N1755, N146);
not NOT1 (N1982, N1968);
and AND4 (N1983, N1978, N1113, N881, N882);
not NOT1 (N1984, N1977);
nand NAND2 (N1985, N1981, N729);
or OR4 (N1986, N1973, N1632, N948, N1278);
xor XOR2 (N1987, N1980, N456);
buf BUF1 (N1988, N1951);
or OR4 (N1989, N1985, N1902, N1018, N1378);
or OR3 (N1990, N1983, N1019, N1099);
or OR3 (N1991, N1982, N135, N1655);
not NOT1 (N1992, N1988);
and AND4 (N1993, N1984, N217, N135, N197);
xor XOR2 (N1994, N1992, N1262);
not NOT1 (N1995, N1965);
or OR3 (N1996, N1993, N1600, N1315);
xor XOR2 (N1997, N1991, N831);
xor XOR2 (N1998, N1996, N530);
or OR2 (N1999, N1994, N110);
not NOT1 (N2000, N1997);
xor XOR2 (N2001, N1987, N525);
not NOT1 (N2002, N1979);
nor NOR3 (N2003, N1989, N1398, N479);
not NOT1 (N2004, N2000);
buf BUF1 (N2005, N2001);
and AND4 (N2006, N1976, N1786, N82, N1958);
buf BUF1 (N2007, N1990);
or OR4 (N2008, N2003, N1476, N706, N531);
or OR4 (N2009, N2005, N1182, N1282, N868);
or OR3 (N2010, N2002, N60, N820);
nand NAND3 (N2011, N2006, N325, N251);
nor NOR3 (N2012, N2011, N1547, N1972);
buf BUF1 (N2013, N2012);
xor XOR2 (N2014, N2010, N1701);
buf BUF1 (N2015, N1999);
buf BUF1 (N2016, N1995);
nand NAND2 (N2017, N2016, N1633);
or OR2 (N2018, N2009, N156);
nor NOR3 (N2019, N2013, N1705, N1318);
xor XOR2 (N2020, N2017, N1808);
xor XOR2 (N2021, N2018, N839);
nor NOR2 (N2022, N1986, N1402);
not NOT1 (N2023, N2021);
buf BUF1 (N2024, N2004);
and AND3 (N2025, N2024, N417, N1834);
and AND4 (N2026, N2020, N1705, N1769, N404);
nor NOR3 (N2027, N2025, N868, N1410);
and AND3 (N2028, N2022, N679, N186);
and AND2 (N2029, N2014, N1720);
nor NOR4 (N2030, N1998, N336, N1724, N795);
xor XOR2 (N2031, N2015, N1078);
nand NAND2 (N2032, N2028, N464);
and AND2 (N2033, N2029, N79);
or OR4 (N2034, N2033, N1201, N1898, N1023);
nor NOR3 (N2035, N2008, N1358, N172);
and AND2 (N2036, N2030, N9);
or OR4 (N2037, N2036, N32, N1736, N539);
and AND2 (N2038, N2032, N740);
buf BUF1 (N2039, N2038);
or OR2 (N2040, N2027, N1632);
buf BUF1 (N2041, N2035);
nand NAND4 (N2042, N2031, N1265, N310, N248);
xor XOR2 (N2043, N2042, N1707);
nor NOR4 (N2044, N2041, N1628, N1334, N1988);
nand NAND4 (N2045, N2044, N1366, N1719, N1869);
xor XOR2 (N2046, N2037, N1152);
or OR2 (N2047, N2026, N1780);
nor NOR3 (N2048, N2047, N80, N1793);
or OR4 (N2049, N2046, N1621, N651, N1578);
nand NAND2 (N2050, N2043, N1735);
not NOT1 (N2051, N2019);
nor NOR3 (N2052, N2048, N1287, N1805);
nand NAND3 (N2053, N2039, N76, N1489);
buf BUF1 (N2054, N2052);
nor NOR3 (N2055, N2054, N1788, N1712);
buf BUF1 (N2056, N2053);
buf BUF1 (N2057, N2049);
nand NAND2 (N2058, N2050, N536);
xor XOR2 (N2059, N2023, N1241);
xor XOR2 (N2060, N2034, N125);
nand NAND3 (N2061, N2045, N66, N561);
and AND2 (N2062, N2059, N615);
nor NOR3 (N2063, N2061, N1976, N131);
and AND4 (N2064, N2062, N571, N1146, N859);
and AND3 (N2065, N2064, N671, N2048);
and AND2 (N2066, N2057, N60);
not NOT1 (N2067, N2051);
or OR3 (N2068, N2056, N1164, N1569);
and AND4 (N2069, N2067, N1487, N1610, N1598);
or OR4 (N2070, N2007, N208, N332, N1963);
nor NOR2 (N2071, N2069, N139);
xor XOR2 (N2072, N2040, N178);
xor XOR2 (N2073, N2070, N1543);
or OR3 (N2074, N2068, N599, N1134);
nand NAND4 (N2075, N2071, N303, N954, N2002);
not NOT1 (N2076, N2065);
nor NOR2 (N2077, N2058, N152);
and AND4 (N2078, N2072, N657, N1802, N2024);
nor NOR4 (N2079, N2077, N149, N1957, N1015);
buf BUF1 (N2080, N2076);
or OR2 (N2081, N2073, N86);
nor NOR3 (N2082, N2055, N2, N573);
and AND2 (N2083, N2066, N426);
nor NOR3 (N2084, N2060, N1860, N230);
buf BUF1 (N2085, N2078);
nand NAND2 (N2086, N2082, N1326);
not NOT1 (N2087, N2085);
nor NOR2 (N2088, N2083, N1623);
buf BUF1 (N2089, N2063);
or OR3 (N2090, N2089, N311, N260);
buf BUF1 (N2091, N2088);
nand NAND2 (N2092, N2080, N710);
buf BUF1 (N2093, N2081);
and AND2 (N2094, N2075, N2020);
and AND4 (N2095, N2086, N232, N742, N1592);
xor XOR2 (N2096, N2092, N196);
nand NAND3 (N2097, N2091, N1110, N1533);
xor XOR2 (N2098, N2090, N1685);
nor NOR4 (N2099, N2097, N235, N215, N801);
xor XOR2 (N2100, N2084, N1297);
nand NAND4 (N2101, N2074, N1572, N499, N710);
xor XOR2 (N2102, N2100, N406);
nand NAND3 (N2103, N2094, N1867, N2064);
xor XOR2 (N2104, N2079, N1342);
nor NOR4 (N2105, N2093, N1520, N468, N1085);
not NOT1 (N2106, N2098);
nand NAND3 (N2107, N2096, N720, N496);
not NOT1 (N2108, N2103);
nand NAND3 (N2109, N2106, N1345, N1656);
xor XOR2 (N2110, N2095, N735);
nand NAND4 (N2111, N2101, N1775, N1459, N1956);
nor NOR2 (N2112, N2110, N393);
nor NOR2 (N2113, N2099, N2006);
nor NOR2 (N2114, N2111, N1391);
nor NOR4 (N2115, N2087, N539, N234, N1756);
and AND4 (N2116, N2113, N2083, N1751, N1805);
nand NAND3 (N2117, N2107, N321, N2089);
nor NOR3 (N2118, N2108, N616, N117);
or OR2 (N2119, N2116, N1341);
not NOT1 (N2120, N2114);
nor NOR4 (N2121, N2112, N1730, N1250, N1316);
nand NAND3 (N2122, N2104, N875, N2089);
not NOT1 (N2123, N2115);
xor XOR2 (N2124, N2118, N1408);
and AND2 (N2125, N2102, N1249);
and AND2 (N2126, N2117, N1019);
not NOT1 (N2127, N2120);
or OR4 (N2128, N2126, N1856, N1624, N2054);
nor NOR4 (N2129, N2125, N1880, N1545, N703);
nand NAND2 (N2130, N2128, N1654);
xor XOR2 (N2131, N2109, N514);
xor XOR2 (N2132, N2123, N572);
and AND3 (N2133, N2122, N1216, N1226);
and AND3 (N2134, N2124, N2096, N975);
nor NOR2 (N2135, N2130, N1249);
and AND2 (N2136, N2135, N346);
or OR2 (N2137, N2121, N1889);
not NOT1 (N2138, N2134);
buf BUF1 (N2139, N2127);
buf BUF1 (N2140, N2129);
nor NOR4 (N2141, N2136, N1091, N1753, N1027);
nand NAND4 (N2142, N2132, N1805, N417, N1598);
buf BUF1 (N2143, N2141);
xor XOR2 (N2144, N2137, N1286);
nand NAND4 (N2145, N2133, N1262, N233, N884);
buf BUF1 (N2146, N2105);
nand NAND4 (N2147, N2138, N839, N1758, N1635);
buf BUF1 (N2148, N2146);
xor XOR2 (N2149, N2119, N1255);
not NOT1 (N2150, N2143);
xor XOR2 (N2151, N2148, N1659);
or OR4 (N2152, N2150, N1594, N853, N955);
nand NAND3 (N2153, N2145, N1727, N1213);
or OR3 (N2154, N2140, N315, N1662);
xor XOR2 (N2155, N2149, N1622);
nor NOR3 (N2156, N2153, N580, N2136);
and AND2 (N2157, N2131, N228);
and AND4 (N2158, N2154, N337, N1002, N624);
nor NOR4 (N2159, N2151, N1084, N1530, N1302);
and AND3 (N2160, N2147, N210, N703);
nor NOR2 (N2161, N2160, N49);
nor NOR2 (N2162, N2161, N1569);
nor NOR3 (N2163, N2142, N887, N1728);
or OR4 (N2164, N2152, N642, N1013, N602);
not NOT1 (N2165, N2158);
and AND3 (N2166, N2155, N717, N1701);
not NOT1 (N2167, N2139);
not NOT1 (N2168, N2163);
or OR2 (N2169, N2164, N1459);
buf BUF1 (N2170, N2162);
and AND2 (N2171, N2157, N812);
or OR2 (N2172, N2171, N141);
buf BUF1 (N2173, N2144);
nor NOR2 (N2174, N2156, N1481);
xor XOR2 (N2175, N2172, N2067);
not NOT1 (N2176, N2170);
or OR3 (N2177, N2168, N2082, N1368);
or OR3 (N2178, N2169, N1471, N652);
and AND2 (N2179, N2176, N1864);
nand NAND2 (N2180, N2166, N532);
buf BUF1 (N2181, N2177);
not NOT1 (N2182, N2173);
buf BUF1 (N2183, N2167);
not NOT1 (N2184, N2180);
not NOT1 (N2185, N2183);
buf BUF1 (N2186, N2185);
buf BUF1 (N2187, N2178);
buf BUF1 (N2188, N2181);
nand NAND4 (N2189, N2184, N895, N1756, N1591);
not NOT1 (N2190, N2174);
or OR4 (N2191, N2189, N1014, N505, N574);
and AND2 (N2192, N2188, N551);
buf BUF1 (N2193, N2182);
nor NOR4 (N2194, N2179, N528, N884, N587);
nor NOR2 (N2195, N2194, N170);
and AND2 (N2196, N2193, N1297);
buf BUF1 (N2197, N2191);
nor NOR4 (N2198, N2192, N1045, N904, N2154);
and AND4 (N2199, N2187, N1108, N952, N201);
nand NAND4 (N2200, N2195, N536, N1339, N1205);
xor XOR2 (N2201, N2197, N225);
not NOT1 (N2202, N2175);
buf BUF1 (N2203, N2202);
xor XOR2 (N2204, N2200, N13);
nor NOR2 (N2205, N2201, N330);
buf BUF1 (N2206, N2199);
not NOT1 (N2207, N2203);
and AND2 (N2208, N2204, N1324);
and AND4 (N2209, N2186, N131, N548, N49);
buf BUF1 (N2210, N2159);
nand NAND4 (N2211, N2165, N1782, N1632, N13);
xor XOR2 (N2212, N2209, N348);
nor NOR4 (N2213, N2196, N405, N670, N1126);
or OR2 (N2214, N2212, N414);
xor XOR2 (N2215, N2198, N2062);
and AND2 (N2216, N2206, N389);
xor XOR2 (N2217, N2211, N1362);
buf BUF1 (N2218, N2214);
not NOT1 (N2219, N2216);
nand NAND4 (N2220, N2213, N1582, N1353, N249);
nor NOR3 (N2221, N2219, N2037, N2021);
xor XOR2 (N2222, N2217, N514);
or OR3 (N2223, N2190, N1927, N1480);
or OR2 (N2224, N2221, N851);
buf BUF1 (N2225, N2223);
not NOT1 (N2226, N2208);
buf BUF1 (N2227, N2215);
not NOT1 (N2228, N2226);
nor NOR3 (N2229, N2222, N427, N243);
not NOT1 (N2230, N2220);
and AND4 (N2231, N2225, N792, N343, N448);
and AND4 (N2232, N2224, N2031, N2155, N2082);
not NOT1 (N2233, N2210);
or OR4 (N2234, N2207, N1464, N765, N1041);
buf BUF1 (N2235, N2228);
buf BUF1 (N2236, N2232);
nor NOR2 (N2237, N2236, N742);
nor NOR4 (N2238, N2227, N1585, N2136, N507);
or OR4 (N2239, N2231, N1834, N113, N393);
buf BUF1 (N2240, N2233);
buf BUF1 (N2241, N2238);
or OR3 (N2242, N2235, N1854, N505);
nand NAND3 (N2243, N2205, N2167, N2136);
not NOT1 (N2244, N2237);
nand NAND3 (N2245, N2234, N1901, N1114);
or OR3 (N2246, N2243, N419, N1533);
and AND4 (N2247, N2239, N1221, N370, N1102);
nor NOR3 (N2248, N2229, N1519, N1603);
or OR3 (N2249, N2247, N1492, N1627);
not NOT1 (N2250, N2245);
xor XOR2 (N2251, N2230, N1719);
xor XOR2 (N2252, N2249, N1811);
and AND2 (N2253, N2241, N1079);
nand NAND2 (N2254, N2253, N1161);
not NOT1 (N2255, N2218);
nand NAND3 (N2256, N2240, N1693, N2129);
nand NAND4 (N2257, N2248, N2114, N804, N322);
buf BUF1 (N2258, N2256);
or OR3 (N2259, N2246, N1999, N544);
nand NAND4 (N2260, N2254, N1632, N1978, N1691);
buf BUF1 (N2261, N2258);
buf BUF1 (N2262, N2252);
not NOT1 (N2263, N2244);
nor NOR4 (N2264, N2257, N1848, N2135, N985);
xor XOR2 (N2265, N2242, N65);
and AND4 (N2266, N2250, N803, N2127, N998);
nor NOR3 (N2267, N2262, N229, N405);
or OR3 (N2268, N2255, N580, N1339);
xor XOR2 (N2269, N2264, N164);
buf BUF1 (N2270, N2268);
or OR2 (N2271, N2263, N661);
nor NOR4 (N2272, N2266, N1969, N1291, N1350);
not NOT1 (N2273, N2251);
nand NAND4 (N2274, N2261, N751, N662, N2051);
nand NAND2 (N2275, N2269, N868);
xor XOR2 (N2276, N2271, N114);
nor NOR4 (N2277, N2272, N2087, N1049, N1752);
nand NAND4 (N2278, N2277, N1185, N392, N1790);
nor NOR3 (N2279, N2276, N1560, N1730);
or OR4 (N2280, N2278, N975, N887, N1708);
and AND4 (N2281, N2274, N1039, N1704, N1045);
nor NOR3 (N2282, N2273, N920, N1925);
xor XOR2 (N2283, N2280, N370);
not NOT1 (N2284, N2260);
buf BUF1 (N2285, N2281);
or OR2 (N2286, N2275, N541);
or OR3 (N2287, N2284, N542, N1782);
nand NAND4 (N2288, N2283, N87, N739, N1826);
not NOT1 (N2289, N2265);
or OR3 (N2290, N2270, N298, N581);
xor XOR2 (N2291, N2290, N1842);
nor NOR3 (N2292, N2285, N852, N1182);
xor XOR2 (N2293, N2282, N1679);
nor NOR3 (N2294, N2289, N1758, N1323);
xor XOR2 (N2295, N2288, N814);
or OR4 (N2296, N2295, N240, N1125, N174);
buf BUF1 (N2297, N2267);
xor XOR2 (N2298, N2292, N491);
xor XOR2 (N2299, N2286, N1864);
xor XOR2 (N2300, N2291, N1849);
xor XOR2 (N2301, N2293, N1889);
buf BUF1 (N2302, N2298);
nor NOR4 (N2303, N2259, N201, N2184, N1219);
nor NOR4 (N2304, N2299, N1430, N1219, N1356);
nand NAND4 (N2305, N2297, N1241, N1621, N349);
xor XOR2 (N2306, N2301, N1550);
buf BUF1 (N2307, N2305);
and AND4 (N2308, N2287, N1566, N9, N264);
not NOT1 (N2309, N2303);
buf BUF1 (N2310, N2309);
nor NOR4 (N2311, N2294, N996, N143, N1537);
nand NAND4 (N2312, N2311, N1738, N426, N1255);
and AND2 (N2313, N2300, N182);
not NOT1 (N2314, N2307);
and AND4 (N2315, N2308, N741, N259, N553);
buf BUF1 (N2316, N2306);
and AND3 (N2317, N2314, N1694, N1737);
and AND3 (N2318, N2315, N772, N1178);
buf BUF1 (N2319, N2312);
and AND4 (N2320, N2279, N964, N871, N602);
and AND2 (N2321, N2318, N2068);
or OR3 (N2322, N2319, N879, N2277);
not NOT1 (N2323, N2302);
not NOT1 (N2324, N2313);
and AND3 (N2325, N2322, N1769, N286);
buf BUF1 (N2326, N2304);
not NOT1 (N2327, N2317);
nand NAND4 (N2328, N2326, N1363, N1048, N1973);
and AND2 (N2329, N2316, N1117);
buf BUF1 (N2330, N2328);
or OR2 (N2331, N2321, N942);
nand NAND2 (N2332, N2310, N1805);
and AND4 (N2333, N2323, N1554, N1608, N1556);
nand NAND4 (N2334, N2330, N1093, N2203, N1975);
buf BUF1 (N2335, N2324);
nor NOR4 (N2336, N2320, N1925, N2065, N1708);
and AND4 (N2337, N2331, N2011, N1306, N818);
nor NOR2 (N2338, N2296, N2076);
not NOT1 (N2339, N2334);
buf BUF1 (N2340, N2339);
or OR3 (N2341, N2338, N1411, N1547);
or OR3 (N2342, N2325, N221, N1692);
not NOT1 (N2343, N2333);
and AND2 (N2344, N2341, N1548);
and AND3 (N2345, N2332, N360, N660);
nor NOR4 (N2346, N2329, N2110, N1307, N2046);
buf BUF1 (N2347, N2340);
buf BUF1 (N2348, N2343);
xor XOR2 (N2349, N2345, N1781);
and AND3 (N2350, N2349, N1118, N1673);
nor NOR3 (N2351, N2344, N2232, N1786);
not NOT1 (N2352, N2347);
nor NOR4 (N2353, N2346, N901, N216, N1343);
xor XOR2 (N2354, N2352, N1888);
nor NOR3 (N2355, N2337, N1132, N440);
nand NAND4 (N2356, N2355, N1869, N649, N1248);
or OR2 (N2357, N2356, N1127);
nand NAND3 (N2358, N2357, N1674, N709);
xor XOR2 (N2359, N2336, N1383);
xor XOR2 (N2360, N2358, N409);
not NOT1 (N2361, N2327);
buf BUF1 (N2362, N2361);
xor XOR2 (N2363, N2342, N1490);
or OR4 (N2364, N2353, N2186, N1289, N2217);
nor NOR4 (N2365, N2348, N839, N679, N1094);
and AND3 (N2366, N2360, N560, N1353);
nor NOR4 (N2367, N2365, N756, N510, N110);
not NOT1 (N2368, N2364);
or OR4 (N2369, N2351, N321, N1776, N193);
not NOT1 (N2370, N2369);
and AND2 (N2371, N2370, N2156);
xor XOR2 (N2372, N2359, N1790);
nand NAND4 (N2373, N2372, N1066, N657, N2088);
and AND3 (N2374, N2367, N1479, N1601);
nand NAND4 (N2375, N2350, N511, N1699, N918);
not NOT1 (N2376, N2363);
and AND3 (N2377, N2362, N982, N2225);
or OR4 (N2378, N2373, N1504, N688, N2008);
not NOT1 (N2379, N2375);
xor XOR2 (N2380, N2376, N1097);
nand NAND2 (N2381, N2378, N756);
nand NAND2 (N2382, N2380, N1898);
not NOT1 (N2383, N2374);
xor XOR2 (N2384, N2368, N2101);
nand NAND3 (N2385, N2366, N2098, N848);
not NOT1 (N2386, N2381);
nand NAND3 (N2387, N2379, N987, N2212);
nor NOR2 (N2388, N2335, N582);
not NOT1 (N2389, N2385);
nor NOR2 (N2390, N2388, N1067);
and AND2 (N2391, N2354, N1289);
buf BUF1 (N2392, N2384);
not NOT1 (N2393, N2392);
buf BUF1 (N2394, N2389);
not NOT1 (N2395, N2387);
not NOT1 (N2396, N2371);
and AND4 (N2397, N2393, N1533, N811, N1945);
xor XOR2 (N2398, N2386, N1088);
xor XOR2 (N2399, N2382, N16);
xor XOR2 (N2400, N2397, N458);
nor NOR3 (N2401, N2391, N236, N2234);
nand NAND3 (N2402, N2394, N1129, N389);
buf BUF1 (N2403, N2400);
and AND3 (N2404, N2377, N65, N175);
buf BUF1 (N2405, N2403);
nor NOR2 (N2406, N2395, N1379);
xor XOR2 (N2407, N2390, N2255);
or OR2 (N2408, N2396, N1126);
or OR4 (N2409, N2401, N2307, N1584, N338);
nor NOR2 (N2410, N2398, N2055);
nor NOR4 (N2411, N2407, N1519, N46, N2207);
buf BUF1 (N2412, N2404);
and AND2 (N2413, N2399, N1302);
nor NOR2 (N2414, N2412, N1688);
or OR2 (N2415, N2406, N622);
xor XOR2 (N2416, N2402, N1902);
nor NOR3 (N2417, N2409, N2197, N1739);
buf BUF1 (N2418, N2383);
nand NAND3 (N2419, N2405, N1749, N499);
not NOT1 (N2420, N2408);
nand NAND4 (N2421, N2413, N1845, N2206, N23);
buf BUF1 (N2422, N2411);
xor XOR2 (N2423, N2420, N1631);
or OR4 (N2424, N2410, N1475, N215, N63);
buf BUF1 (N2425, N2417);
or OR4 (N2426, N2414, N1976, N1375, N843);
and AND3 (N2427, N2425, N1715, N429);
not NOT1 (N2428, N2415);
nand NAND3 (N2429, N2422, N155, N1106);
xor XOR2 (N2430, N2429, N1150);
buf BUF1 (N2431, N2424);
and AND2 (N2432, N2431, N150);
not NOT1 (N2433, N2423);
nand NAND4 (N2434, N2426, N338, N1309, N1694);
buf BUF1 (N2435, N2433);
nand NAND2 (N2436, N2435, N2427);
or OR4 (N2437, N634, N1618, N967, N1698);
xor XOR2 (N2438, N2436, N548);
nand NAND4 (N2439, N2428, N1729, N378, N1727);
nor NOR4 (N2440, N2430, N2002, N2001, N155);
and AND4 (N2441, N2432, N1500, N489, N1384);
nand NAND2 (N2442, N2441, N134);
and AND3 (N2443, N2419, N1027, N1761);
nor NOR2 (N2444, N2418, N2140);
buf BUF1 (N2445, N2444);
nor NOR2 (N2446, N2440, N765);
xor XOR2 (N2447, N2421, N1422);
buf BUF1 (N2448, N2447);
nand NAND2 (N2449, N2448, N2200);
nor NOR3 (N2450, N2445, N1889, N2217);
nor NOR2 (N2451, N2446, N1896);
xor XOR2 (N2452, N2416, N1364);
or OR3 (N2453, N2442, N857, N1571);
or OR2 (N2454, N2449, N1284);
nand NAND2 (N2455, N2434, N2088);
not NOT1 (N2456, N2451);
buf BUF1 (N2457, N2456);
buf BUF1 (N2458, N2455);
nor NOR4 (N2459, N2457, N599, N2018, N1054);
nor NOR3 (N2460, N2452, N873, N1304);
xor XOR2 (N2461, N2450, N2106);
nand NAND3 (N2462, N2454, N1949, N1782);
or OR3 (N2463, N2438, N907, N1746);
buf BUF1 (N2464, N2453);
and AND3 (N2465, N2458, N1362, N1211);
or OR3 (N2466, N2439, N366, N1150);
or OR3 (N2467, N2437, N1226, N1109);
and AND3 (N2468, N2467, N1880, N41);
xor XOR2 (N2469, N2468, N1330);
not NOT1 (N2470, N2464);
nor NOR2 (N2471, N2465, N1610);
buf BUF1 (N2472, N2471);
or OR3 (N2473, N2461, N1675, N2333);
nand NAND2 (N2474, N2469, N712);
not NOT1 (N2475, N2443);
or OR3 (N2476, N2459, N1652, N1543);
nand NAND2 (N2477, N2470, N1594);
nand NAND2 (N2478, N2466, N2413);
xor XOR2 (N2479, N2462, N1074);
and AND3 (N2480, N2472, N750, N2221);
xor XOR2 (N2481, N2477, N2314);
nor NOR3 (N2482, N2463, N512, N1713);
nor NOR4 (N2483, N2475, N8, N2037, N1269);
nor NOR4 (N2484, N2473, N1337, N1229, N391);
not NOT1 (N2485, N2476);
nand NAND4 (N2486, N2485, N596, N798, N1532);
nor NOR4 (N2487, N2484, N1089, N474, N86);
and AND3 (N2488, N2481, N1042, N970);
nor NOR3 (N2489, N2474, N122, N1974);
nor NOR4 (N2490, N2487, N1552, N1817, N2014);
or OR2 (N2491, N2482, N2054);
xor XOR2 (N2492, N2460, N180);
buf BUF1 (N2493, N2491);
and AND4 (N2494, N2480, N2229, N170, N1852);
buf BUF1 (N2495, N2494);
not NOT1 (N2496, N2495);
nand NAND4 (N2497, N2490, N2072, N657, N347);
or OR3 (N2498, N2492, N582, N1758);
nor NOR2 (N2499, N2489, N1695);
buf BUF1 (N2500, N2493);
xor XOR2 (N2501, N2486, N1183);
xor XOR2 (N2502, N2498, N497);
and AND2 (N2503, N2496, N2310);
not NOT1 (N2504, N2503);
buf BUF1 (N2505, N2497);
not NOT1 (N2506, N2505);
buf BUF1 (N2507, N2478);
and AND4 (N2508, N2500, N29, N921, N784);
nor NOR4 (N2509, N2507, N840, N751, N138);
not NOT1 (N2510, N2509);
buf BUF1 (N2511, N2488);
or OR3 (N2512, N2499, N1975, N1321);
or OR4 (N2513, N2502, N1037, N85, N291);
xor XOR2 (N2514, N2504, N1527);
not NOT1 (N2515, N2511);
nor NOR4 (N2516, N2515, N1825, N459, N1741);
nand NAND4 (N2517, N2501, N1397, N1434, N408);
and AND4 (N2518, N2483, N2356, N1123, N837);
xor XOR2 (N2519, N2510, N589);
xor XOR2 (N2520, N2479, N1239);
buf BUF1 (N2521, N2520);
buf BUF1 (N2522, N2512);
not NOT1 (N2523, N2519);
or OR3 (N2524, N2521, N1988, N1186);
nor NOR4 (N2525, N2523, N2229, N355, N701);
xor XOR2 (N2526, N2506, N321);
nand NAND4 (N2527, N2518, N1229, N93, N1021);
buf BUF1 (N2528, N2525);
or OR3 (N2529, N2508, N2267, N1695);
nor NOR3 (N2530, N2529, N2071, N1530);
or OR4 (N2531, N2516, N1435, N1464, N1973);
nand NAND3 (N2532, N2524, N2176, N146);
nor NOR4 (N2533, N2517, N2195, N2336, N1725);
xor XOR2 (N2534, N2528, N764);
or OR3 (N2535, N2526, N1612, N178);
not NOT1 (N2536, N2535);
buf BUF1 (N2537, N2530);
nand NAND2 (N2538, N2514, N1175);
nand NAND4 (N2539, N2522, N19, N2202, N1956);
nor NOR3 (N2540, N2531, N1867, N1481);
nor NOR3 (N2541, N2538, N636, N396);
or OR2 (N2542, N2513, N1670);
or OR3 (N2543, N2533, N2541, N921);
buf BUF1 (N2544, N1582);
nor NOR3 (N2545, N2543, N1892, N1470);
xor XOR2 (N2546, N2536, N121);
and AND2 (N2547, N2544, N1095);
and AND4 (N2548, N2532, N1903, N394, N1787);
or OR3 (N2549, N2527, N507, N822);
or OR4 (N2550, N2537, N166, N1026, N54);
xor XOR2 (N2551, N2539, N1551);
and AND2 (N2552, N2547, N2405);
nor NOR4 (N2553, N2551, N564, N268, N1492);
nand NAND2 (N2554, N2542, N515);
xor XOR2 (N2555, N2546, N877);
or OR2 (N2556, N2548, N79);
or OR4 (N2557, N2549, N1452, N2166, N929);
or OR4 (N2558, N2553, N88, N156, N642);
or OR3 (N2559, N2558, N878, N469);
buf BUF1 (N2560, N2540);
or OR3 (N2561, N2550, N527, N699);
nor NOR4 (N2562, N2557, N1684, N816, N2426);
nor NOR3 (N2563, N2554, N2170, N731);
nor NOR3 (N2564, N2534, N1813, N804);
or OR4 (N2565, N2556, N1926, N2001, N213);
xor XOR2 (N2566, N2560, N1163);
nor NOR4 (N2567, N2562, N2170, N1997, N559);
or OR3 (N2568, N2563, N468, N2507);
or OR4 (N2569, N2555, N2355, N1470, N364);
xor XOR2 (N2570, N2564, N934);
xor XOR2 (N2571, N2568, N2077);
nor NOR4 (N2572, N2569, N339, N470, N297);
and AND2 (N2573, N2565, N2509);
buf BUF1 (N2574, N2561);
not NOT1 (N2575, N2572);
and AND2 (N2576, N2570, N338);
xor XOR2 (N2577, N2566, N2047);
nand NAND2 (N2578, N2559, N754);
buf BUF1 (N2579, N2578);
or OR3 (N2580, N2577, N2259, N436);
nand NAND3 (N2581, N2573, N2398, N607);
buf BUF1 (N2582, N2579);
not NOT1 (N2583, N2575);
buf BUF1 (N2584, N2581);
not NOT1 (N2585, N2580);
nor NOR2 (N2586, N2567, N1408);
and AND2 (N2587, N2545, N96);
buf BUF1 (N2588, N2571);
and AND2 (N2589, N2576, N500);
not NOT1 (N2590, N2587);
buf BUF1 (N2591, N2552);
buf BUF1 (N2592, N2574);
and AND4 (N2593, N2588, N1200, N1184, N2286);
not NOT1 (N2594, N2590);
nand NAND2 (N2595, N2584, N1920);
buf BUF1 (N2596, N2585);
or OR3 (N2597, N2591, N1729, N140);
and AND4 (N2598, N2594, N2254, N809, N2587);
nor NOR4 (N2599, N2593, N446, N1269, N2236);
nor NOR3 (N2600, N2592, N1839, N637);
buf BUF1 (N2601, N2586);
or OR4 (N2602, N2599, N871, N558, N2308);
buf BUF1 (N2603, N2602);
xor XOR2 (N2604, N2596, N2490);
not NOT1 (N2605, N2603);
and AND2 (N2606, N2595, N1642);
not NOT1 (N2607, N2605);
or OR3 (N2608, N2597, N1864, N715);
xor XOR2 (N2609, N2598, N151);
buf BUF1 (N2610, N2609);
not NOT1 (N2611, N2589);
nor NOR3 (N2612, N2600, N1967, N990);
or OR2 (N2613, N2582, N2565);
or OR3 (N2614, N2612, N1925, N1851);
or OR2 (N2615, N2583, N108);
buf BUF1 (N2616, N2614);
xor XOR2 (N2617, N2604, N2423);
xor XOR2 (N2618, N2607, N817);
xor XOR2 (N2619, N2618, N1332);
not NOT1 (N2620, N2601);
and AND2 (N2621, N2617, N2489);
nor NOR3 (N2622, N2606, N2048, N777);
and AND4 (N2623, N2619, N117, N1786, N2257);
xor XOR2 (N2624, N2616, N1934);
and AND3 (N2625, N2620, N208, N1781);
or OR2 (N2626, N2625, N764);
and AND2 (N2627, N2623, N2570);
nor NOR4 (N2628, N2611, N2581, N1597, N2183);
not NOT1 (N2629, N2621);
and AND2 (N2630, N2626, N1197);
and AND2 (N2631, N2608, N774);
not NOT1 (N2632, N2628);
xor XOR2 (N2633, N2615, N1070);
and AND3 (N2634, N2631, N325, N1122);
and AND2 (N2635, N2629, N1453);
and AND4 (N2636, N2613, N1402, N666, N2617);
nor NOR4 (N2637, N2622, N2173, N2182, N680);
buf BUF1 (N2638, N2635);
xor XOR2 (N2639, N2634, N1565);
xor XOR2 (N2640, N2633, N1806);
or OR2 (N2641, N2637, N1266);
xor XOR2 (N2642, N2636, N1286);
not NOT1 (N2643, N2642);
not NOT1 (N2644, N2641);
nand NAND4 (N2645, N2640, N504, N2317, N536);
not NOT1 (N2646, N2632);
and AND3 (N2647, N2645, N883, N1209);
nand NAND4 (N2648, N2643, N1178, N633, N852);
nand NAND2 (N2649, N2627, N2339);
buf BUF1 (N2650, N2610);
not NOT1 (N2651, N2624);
and AND3 (N2652, N2647, N2442, N1892);
xor XOR2 (N2653, N2646, N1415);
nor NOR3 (N2654, N2639, N1798, N183);
and AND4 (N2655, N2651, N1708, N387, N307);
nor NOR3 (N2656, N2655, N1732, N1213);
nor NOR2 (N2657, N2654, N2091);
or OR3 (N2658, N2648, N2269, N2278);
buf BUF1 (N2659, N2650);
or OR3 (N2660, N2630, N1502, N524);
buf BUF1 (N2661, N2652);
xor XOR2 (N2662, N2638, N2619);
xor XOR2 (N2663, N2644, N1146);
not NOT1 (N2664, N2663);
buf BUF1 (N2665, N2662);
nor NOR2 (N2666, N2649, N126);
not NOT1 (N2667, N2659);
nand NAND2 (N2668, N2657, N2143);
not NOT1 (N2669, N2668);
nor NOR4 (N2670, N2653, N972, N130, N787);
and AND2 (N2671, N2667, N2038);
xor XOR2 (N2672, N2661, N1118);
nand NAND3 (N2673, N2671, N1941, N1561);
and AND4 (N2674, N2658, N1331, N760, N2658);
buf BUF1 (N2675, N2660);
xor XOR2 (N2676, N2669, N1191);
xor XOR2 (N2677, N2656, N108);
nand NAND4 (N2678, N2666, N1462, N1248, N141);
not NOT1 (N2679, N2665);
buf BUF1 (N2680, N2675);
xor XOR2 (N2681, N2680, N2068);
buf BUF1 (N2682, N2672);
xor XOR2 (N2683, N2676, N1833);
not NOT1 (N2684, N2682);
and AND3 (N2685, N2679, N1110, N1824);
xor XOR2 (N2686, N2678, N375);
nand NAND3 (N2687, N2664, N2211, N707);
not NOT1 (N2688, N2683);
nand NAND3 (N2689, N2677, N864, N2375);
or OR2 (N2690, N2684, N2540);
or OR2 (N2691, N2689, N1362);
nand NAND2 (N2692, N2690, N2055);
buf BUF1 (N2693, N2685);
nor NOR4 (N2694, N2693, N155, N478, N1990);
or OR2 (N2695, N2694, N927);
or OR3 (N2696, N2691, N1366, N2221);
or OR3 (N2697, N2670, N1816, N1168);
and AND4 (N2698, N2673, N1694, N184, N1373);
nor NOR3 (N2699, N2674, N1690, N2003);
buf BUF1 (N2700, N2692);
nor NOR3 (N2701, N2688, N1927, N471);
xor XOR2 (N2702, N2699, N2577);
not NOT1 (N2703, N2697);
or OR3 (N2704, N2681, N11, N734);
buf BUF1 (N2705, N2703);
and AND2 (N2706, N2687, N1416);
xor XOR2 (N2707, N2686, N2374);
nand NAND3 (N2708, N2705, N1648, N449);
nor NOR3 (N2709, N2695, N2415, N428);
not NOT1 (N2710, N2708);
nor NOR4 (N2711, N2706, N1349, N581, N250);
xor XOR2 (N2712, N2711, N253);
nor NOR3 (N2713, N2698, N371, N1994);
or OR2 (N2714, N2710, N1199);
nor NOR3 (N2715, N2707, N1355, N1764);
and AND2 (N2716, N2713, N8);
nor NOR4 (N2717, N2696, N750, N2376, N2673);
nor NOR4 (N2718, N2701, N2370, N2247, N2074);
nor NOR4 (N2719, N2704, N2323, N711, N412);
nand NAND2 (N2720, N2717, N111);
or OR3 (N2721, N2715, N2131, N2335);
not NOT1 (N2722, N2718);
not NOT1 (N2723, N2720);
xor XOR2 (N2724, N2716, N1415);
nor NOR3 (N2725, N2709, N369, N933);
nand NAND3 (N2726, N2724, N2523, N83);
not NOT1 (N2727, N2722);
xor XOR2 (N2728, N2719, N1278);
nor NOR3 (N2729, N2728, N2667, N1634);
not NOT1 (N2730, N2721);
nand NAND3 (N2731, N2726, N2578, N1905);
nor NOR3 (N2732, N2731, N346, N1762);
nor NOR2 (N2733, N2732, N71);
xor XOR2 (N2734, N2727, N2006);
and AND4 (N2735, N2723, N449, N674, N308);
nand NAND3 (N2736, N2733, N211, N467);
nand NAND3 (N2737, N2725, N909, N2654);
nand NAND3 (N2738, N2734, N1371, N1628);
xor XOR2 (N2739, N2729, N41);
and AND2 (N2740, N2738, N1486);
nor NOR4 (N2741, N2740, N2560, N2143, N223);
or OR2 (N2742, N2737, N1208);
or OR3 (N2743, N2730, N1232, N2627);
xor XOR2 (N2744, N2735, N62);
xor XOR2 (N2745, N2743, N2371);
nand NAND3 (N2746, N2744, N784, N457);
xor XOR2 (N2747, N2742, N1933);
and AND4 (N2748, N2714, N2320, N76, N2686);
and AND2 (N2749, N2712, N1519);
and AND4 (N2750, N2739, N167, N968, N668);
or OR4 (N2751, N2741, N2576, N2685, N1671);
buf BUF1 (N2752, N2700);
and AND2 (N2753, N2750, N553);
nor NOR3 (N2754, N2746, N508, N539);
or OR4 (N2755, N2745, N465, N2661, N1651);
xor XOR2 (N2756, N2749, N2202);
nor NOR4 (N2757, N2753, N127, N1449, N786);
not NOT1 (N2758, N2754);
buf BUF1 (N2759, N2747);
xor XOR2 (N2760, N2758, N2537);
and AND2 (N2761, N2752, N445);
xor XOR2 (N2762, N2702, N2628);
xor XOR2 (N2763, N2755, N1448);
buf BUF1 (N2764, N2736);
buf BUF1 (N2765, N2756);
or OR2 (N2766, N2761, N2217);
nand NAND2 (N2767, N2766, N1792);
or OR4 (N2768, N2767, N2061, N521, N1918);
nor NOR4 (N2769, N2757, N2026, N357, N1441);
nand NAND3 (N2770, N2764, N1479, N2092);
and AND2 (N2771, N2768, N1026);
buf BUF1 (N2772, N2770);
nand NAND2 (N2773, N2772, N1443);
nor NOR4 (N2774, N2751, N4, N1321, N965);
nand NAND2 (N2775, N2762, N2598);
and AND3 (N2776, N2775, N1139, N1753);
buf BUF1 (N2777, N2774);
buf BUF1 (N2778, N2748);
not NOT1 (N2779, N2777);
buf BUF1 (N2780, N2759);
nor NOR4 (N2781, N2778, N654, N105, N853);
nor NOR3 (N2782, N2765, N2636, N97);
or OR4 (N2783, N2773, N115, N1304, N2543);
not NOT1 (N2784, N2763);
nand NAND3 (N2785, N2779, N475, N328);
xor XOR2 (N2786, N2776, N2206);
buf BUF1 (N2787, N2783);
or OR2 (N2788, N2769, N1903);
or OR2 (N2789, N2781, N598);
xor XOR2 (N2790, N2784, N1165);
xor XOR2 (N2791, N2788, N961);
buf BUF1 (N2792, N2782);
nor NOR3 (N2793, N2760, N2631, N2042);
buf BUF1 (N2794, N2786);
and AND3 (N2795, N2771, N448, N2321);
nand NAND2 (N2796, N2794, N990);
buf BUF1 (N2797, N2789);
not NOT1 (N2798, N2796);
buf BUF1 (N2799, N2780);
xor XOR2 (N2800, N2795, N1178);
buf BUF1 (N2801, N2793);
nand NAND3 (N2802, N2787, N1647, N1398);
xor XOR2 (N2803, N2797, N255);
and AND4 (N2804, N2798, N2422, N2018, N1305);
nand NAND2 (N2805, N2791, N1189);
nand NAND3 (N2806, N2803, N2037, N2415);
or OR4 (N2807, N2790, N1820, N1134, N1387);
nand NAND4 (N2808, N2800, N452, N1209, N1920);
xor XOR2 (N2809, N2785, N309);
nand NAND2 (N2810, N2802, N93);
not NOT1 (N2811, N2801);
nand NAND4 (N2812, N2792, N396, N533, N2245);
or OR4 (N2813, N2804, N453, N599, N96);
not NOT1 (N2814, N2805);
not NOT1 (N2815, N2807);
not NOT1 (N2816, N2810);
nand NAND3 (N2817, N2813, N1907, N135);
or OR4 (N2818, N2812, N753, N283, N2465);
buf BUF1 (N2819, N2799);
not NOT1 (N2820, N2818);
xor XOR2 (N2821, N2815, N808);
xor XOR2 (N2822, N2821, N408);
or OR2 (N2823, N2820, N30);
xor XOR2 (N2824, N2808, N1684);
nor NOR2 (N2825, N2824, N136);
buf BUF1 (N2826, N2816);
nand NAND4 (N2827, N2825, N120, N1655, N1750);
nor NOR3 (N2828, N2809, N1095, N1162);
not NOT1 (N2829, N2828);
nand NAND3 (N2830, N2819, N2653, N2351);
not NOT1 (N2831, N2811);
nand NAND4 (N2832, N2829, N2138, N2033, N288);
not NOT1 (N2833, N2826);
or OR2 (N2834, N2831, N823);
not NOT1 (N2835, N2833);
buf BUF1 (N2836, N2830);
nand NAND4 (N2837, N2827, N2095, N1922, N1310);
not NOT1 (N2838, N2822);
nor NOR3 (N2839, N2838, N114, N1177);
not NOT1 (N2840, N2835);
xor XOR2 (N2841, N2832, N759);
or OR2 (N2842, N2841, N160);
or OR4 (N2843, N2842, N379, N602, N1254);
nand NAND2 (N2844, N2843, N477);
nand NAND4 (N2845, N2844, N2351, N844, N2504);
nor NOR2 (N2846, N2817, N562);
or OR4 (N2847, N2839, N760, N188, N2463);
buf BUF1 (N2848, N2836);
and AND2 (N2849, N2848, N231);
nor NOR3 (N2850, N2849, N739, N1656);
nor NOR4 (N2851, N2840, N1160, N2374, N655);
not NOT1 (N2852, N2846);
nor NOR3 (N2853, N2845, N2304, N2082);
and AND4 (N2854, N2853, N752, N717, N262);
or OR3 (N2855, N2814, N2328, N170);
nor NOR2 (N2856, N2806, N2511);
buf BUF1 (N2857, N2823);
not NOT1 (N2858, N2852);
xor XOR2 (N2859, N2855, N750);
nand NAND3 (N2860, N2858, N1051, N1278);
or OR4 (N2861, N2859, N1639, N2625, N1514);
buf BUF1 (N2862, N2850);
and AND4 (N2863, N2834, N1442, N2249, N2593);
nor NOR4 (N2864, N2837, N1756, N1215, N846);
and AND4 (N2865, N2860, N757, N341, N537);
not NOT1 (N2866, N2847);
or OR3 (N2867, N2864, N2050, N2653);
xor XOR2 (N2868, N2863, N578);
or OR2 (N2869, N2857, N791);
or OR3 (N2870, N2865, N2545, N477);
not NOT1 (N2871, N2851);
or OR4 (N2872, N2861, N2203, N1712, N1004);
nand NAND3 (N2873, N2870, N737, N428);
or OR3 (N2874, N2867, N2845, N1108);
xor XOR2 (N2875, N2869, N1140);
nand NAND3 (N2876, N2875, N2587, N460);
or OR3 (N2877, N2873, N911, N700);
buf BUF1 (N2878, N2871);
and AND3 (N2879, N2877, N1572, N1108);
not NOT1 (N2880, N2866);
xor XOR2 (N2881, N2856, N1459);
or OR3 (N2882, N2878, N1937, N1064);
or OR2 (N2883, N2862, N1930);
and AND4 (N2884, N2879, N2594, N2298, N2137);
buf BUF1 (N2885, N2854);
nor NOR4 (N2886, N2882, N613, N1768, N2575);
or OR3 (N2887, N2884, N2096, N1364);
not NOT1 (N2888, N2872);
buf BUF1 (N2889, N2876);
nor NOR3 (N2890, N2888, N1813, N577);
or OR3 (N2891, N2887, N2812, N1087);
and AND2 (N2892, N2885, N1962);
and AND4 (N2893, N2874, N84, N578, N2645);
not NOT1 (N2894, N2893);
buf BUF1 (N2895, N2883);
xor XOR2 (N2896, N2891, N641);
buf BUF1 (N2897, N2890);
xor XOR2 (N2898, N2896, N172);
nor NOR2 (N2899, N2868, N1457);
not NOT1 (N2900, N2899);
nand NAND4 (N2901, N2895, N2538, N2317, N1047);
nand NAND4 (N2902, N2898, N808, N1913, N1897);
or OR2 (N2903, N2901, N1084);
not NOT1 (N2904, N2881);
not NOT1 (N2905, N2886);
xor XOR2 (N2906, N2900, N2061);
nor NOR2 (N2907, N2894, N2287);
nor NOR3 (N2908, N2905, N1637, N717);
nand NAND4 (N2909, N2907, N1362, N2606, N262);
and AND4 (N2910, N2908, N379, N2610, N291);
nand NAND3 (N2911, N2892, N2687, N2317);
or OR2 (N2912, N2904, N588);
buf BUF1 (N2913, N2911);
buf BUF1 (N2914, N2903);
buf BUF1 (N2915, N2880);
or OR3 (N2916, N2913, N103, N2612);
nor NOR3 (N2917, N2915, N180, N1659);
or OR2 (N2918, N2897, N1751);
xor XOR2 (N2919, N2889, N2686);
or OR4 (N2920, N2914, N1825, N1565, N1465);
and AND3 (N2921, N2909, N2175, N680);
nor NOR3 (N2922, N2917, N1630, N2184);
and AND4 (N2923, N2902, N2134, N1151, N498);
not NOT1 (N2924, N2906);
nor NOR2 (N2925, N2920, N1915);
nor NOR3 (N2926, N2912, N1103, N1827);
nor NOR3 (N2927, N2918, N1449, N2564);
nand NAND3 (N2928, N2919, N545, N2212);
nor NOR3 (N2929, N2916, N2174, N2194);
nor NOR4 (N2930, N2929, N2308, N460, N350);
not NOT1 (N2931, N2928);
or OR2 (N2932, N2931, N1098);
or OR3 (N2933, N2924, N1014, N1398);
xor XOR2 (N2934, N2925, N2331);
or OR2 (N2935, N2922, N15);
and AND4 (N2936, N2910, N24, N623, N1618);
buf BUF1 (N2937, N2932);
and AND4 (N2938, N2927, N784, N2716, N1458);
or OR4 (N2939, N2938, N115, N2898, N1157);
nor NOR4 (N2940, N2934, N293, N1290, N1939);
not NOT1 (N2941, N2933);
nand NAND2 (N2942, N2930, N1232);
not NOT1 (N2943, N2921);
nand NAND3 (N2944, N2926, N1757, N145);
nand NAND3 (N2945, N2944, N2194, N1256);
or OR2 (N2946, N2937, N2426);
nor NOR3 (N2947, N2943, N737, N210);
nand NAND4 (N2948, N2941, N685, N32, N1356);
and AND4 (N2949, N2942, N900, N1755, N2434);
or OR2 (N2950, N2945, N1531);
xor XOR2 (N2951, N2923, N1911);
or OR4 (N2952, N2948, N1979, N1419, N486);
not NOT1 (N2953, N2935);
or OR3 (N2954, N2936, N1891, N1684);
not NOT1 (N2955, N2940);
buf BUF1 (N2956, N2947);
nor NOR4 (N2957, N2956, N1360, N632, N2543);
not NOT1 (N2958, N2946);
buf BUF1 (N2959, N2953);
xor XOR2 (N2960, N2949, N2778);
xor XOR2 (N2961, N2960, N2286);
xor XOR2 (N2962, N2939, N2667);
not NOT1 (N2963, N2962);
buf BUF1 (N2964, N2959);
not NOT1 (N2965, N2952);
buf BUF1 (N2966, N2954);
nand NAND4 (N2967, N2950, N754, N281, N1640);
not NOT1 (N2968, N2964);
and AND4 (N2969, N2968, N750, N1100, N47);
nand NAND2 (N2970, N2955, N27);
or OR2 (N2971, N2965, N1056);
nor NOR3 (N2972, N2969, N2745, N1008);
or OR3 (N2973, N2971, N1156, N495);
nand NAND2 (N2974, N2963, N2416);
or OR3 (N2975, N2958, N1745, N1563);
nor NOR3 (N2976, N2966, N1538, N1893);
xor XOR2 (N2977, N2970, N512);
nand NAND4 (N2978, N2975, N2069, N566, N301);
nand NAND3 (N2979, N2957, N922, N1539);
not NOT1 (N2980, N2979);
and AND2 (N2981, N2951, N2959);
not NOT1 (N2982, N2978);
nor NOR4 (N2983, N2977, N1260, N2056, N444);
buf BUF1 (N2984, N2982);
or OR2 (N2985, N2972, N1953);
buf BUF1 (N2986, N2967);
nor NOR4 (N2987, N2983, N103, N2162, N2479);
nand NAND4 (N2988, N2984, N702, N1835, N1014);
xor XOR2 (N2989, N2973, N650);
or OR2 (N2990, N2986, N2287);
xor XOR2 (N2991, N2981, N1552);
or OR3 (N2992, N2980, N1542, N1341);
not NOT1 (N2993, N2992);
xor XOR2 (N2994, N2976, N61);
nand NAND4 (N2995, N2993, N92, N160, N1357);
and AND4 (N2996, N2987, N1937, N1201, N190);
nand NAND2 (N2997, N2961, N1429);
and AND2 (N2998, N2994, N1407);
or OR2 (N2999, N2997, N1365);
xor XOR2 (N3000, N2989, N932);
or OR3 (N3001, N2998, N2431, N2651);
nor NOR4 (N3002, N3000, N978, N2262, N1560);
and AND4 (N3003, N2974, N1376, N2847, N2192);
buf BUF1 (N3004, N2999);
nand NAND3 (N3005, N2995, N805, N2705);
nand NAND4 (N3006, N3004, N722, N278, N2704);
xor XOR2 (N3007, N3003, N1261);
or OR4 (N3008, N3005, N290, N1460, N1415);
and AND4 (N3009, N3006, N1206, N858, N1459);
nand NAND4 (N3010, N3002, N1725, N1554, N1430);
or OR4 (N3011, N2988, N2404, N319, N947);
and AND4 (N3012, N2985, N482, N1593, N2101);
xor XOR2 (N3013, N3008, N1168);
or OR3 (N3014, N3009, N1494, N986);
nor NOR4 (N3015, N3010, N1711, N1127, N2639);
xor XOR2 (N3016, N2990, N2550);
nor NOR4 (N3017, N3001, N1793, N1726, N2113);
and AND2 (N3018, N3007, N227);
buf BUF1 (N3019, N3017);
buf BUF1 (N3020, N3014);
or OR3 (N3021, N3019, N476, N1790);
xor XOR2 (N3022, N3015, N1576);
nor NOR4 (N3023, N3011, N1987, N1937, N917);
or OR2 (N3024, N3012, N2530);
nand NAND4 (N3025, N3018, N2573, N1053, N1640);
and AND2 (N3026, N3025, N1812);
xor XOR2 (N3027, N3020, N1566);
nor NOR2 (N3028, N3022, N1320);
and AND4 (N3029, N3023, N559, N343, N913);
not NOT1 (N3030, N3029);
nand NAND2 (N3031, N3013, N1526);
nor NOR4 (N3032, N3021, N2078, N462, N1504);
nor NOR4 (N3033, N3027, N313, N1695, N88);
and AND2 (N3034, N3028, N2176);
and AND2 (N3035, N3033, N171);
or OR2 (N3036, N3034, N1125);
not NOT1 (N3037, N3031);
not NOT1 (N3038, N3030);
not NOT1 (N3039, N3032);
xor XOR2 (N3040, N3035, N2668);
nor NOR4 (N3041, N2996, N34, N2083, N1639);
nor NOR4 (N3042, N3041, N1474, N2434, N820);
nand NAND3 (N3043, N3042, N1010, N3019);
nand NAND4 (N3044, N3039, N2935, N2555, N1372);
not NOT1 (N3045, N2991);
nor NOR3 (N3046, N3016, N1298, N2650);
buf BUF1 (N3047, N3038);
and AND4 (N3048, N3044, N2352, N2406, N1222);
and AND4 (N3049, N3047, N2275, N554, N2239);
and AND4 (N3050, N3026, N522, N1635, N2978);
nor NOR4 (N3051, N3045, N697, N2432, N1539);
nand NAND2 (N3052, N3037, N1957);
buf BUF1 (N3053, N3040);
nor NOR3 (N3054, N3053, N1472, N2893);
not NOT1 (N3055, N3048);
xor XOR2 (N3056, N3051, N2658);
nand NAND4 (N3057, N3043, N1704, N482, N749);
and AND2 (N3058, N3055, N2286);
nor NOR2 (N3059, N3046, N1538);
or OR4 (N3060, N3024, N1529, N701, N683);
buf BUF1 (N3061, N3036);
and AND4 (N3062, N3058, N1712, N488, N1984);
buf BUF1 (N3063, N3059);
buf BUF1 (N3064, N3061);
and AND4 (N3065, N3050, N2836, N68, N493);
and AND3 (N3066, N3057, N716, N83);
and AND2 (N3067, N3065, N1857);
xor XOR2 (N3068, N3063, N1480);
not NOT1 (N3069, N3068);
xor XOR2 (N3070, N3060, N690);
buf BUF1 (N3071, N3049);
or OR4 (N3072, N3070, N2336, N956, N465);
nor NOR3 (N3073, N3071, N910, N91);
not NOT1 (N3074, N3073);
nor NOR3 (N3075, N3062, N1126, N2597);
not NOT1 (N3076, N3054);
not NOT1 (N3077, N3076);
not NOT1 (N3078, N3066);
xor XOR2 (N3079, N3075, N1170);
xor XOR2 (N3080, N3077, N2069);
not NOT1 (N3081, N3064);
nand NAND4 (N3082, N3072, N1095, N738, N1765);
and AND3 (N3083, N3081, N1239, N1120);
nand NAND3 (N3084, N3083, N742, N2489);
or OR4 (N3085, N3052, N2307, N2388, N2665);
and AND2 (N3086, N3082, N901);
or OR4 (N3087, N3074, N814, N2939, N2251);
or OR3 (N3088, N3086, N1096, N418);
or OR3 (N3089, N3067, N2818, N1484);
and AND4 (N3090, N3087, N883, N1348, N327);
xor XOR2 (N3091, N3088, N579);
xor XOR2 (N3092, N3089, N2842);
or OR2 (N3093, N3078, N1939);
xor XOR2 (N3094, N3093, N1613);
or OR4 (N3095, N3084, N14, N2653, N2036);
nand NAND3 (N3096, N3080, N1862, N2512);
or OR3 (N3097, N3092, N651, N1833);
or OR4 (N3098, N3095, N877, N582, N1598);
nand NAND2 (N3099, N3069, N743);
buf BUF1 (N3100, N3099);
nor NOR4 (N3101, N3098, N1978, N1478, N42);
xor XOR2 (N3102, N3091, N2421);
buf BUF1 (N3103, N3094);
nor NOR2 (N3104, N3102, N1939);
nand NAND4 (N3105, N3104, N182, N805, N2176);
nand NAND2 (N3106, N3105, N958);
buf BUF1 (N3107, N3100);
not NOT1 (N3108, N3097);
or OR4 (N3109, N3108, N2242, N98, N3030);
xor XOR2 (N3110, N3109, N1722);
nor NOR2 (N3111, N3110, N2377);
or OR4 (N3112, N3107, N1465, N2137, N1536);
buf BUF1 (N3113, N3085);
and AND2 (N3114, N3101, N979);
and AND3 (N3115, N3112, N2919, N631);
or OR4 (N3116, N3079, N460, N2283, N2727);
buf BUF1 (N3117, N3115);
nor NOR2 (N3118, N3096, N1738);
and AND2 (N3119, N3103, N172);
nand NAND2 (N3120, N3056, N1563);
nand NAND3 (N3121, N3120, N345, N1520);
and AND3 (N3122, N3111, N258, N1492);
or OR2 (N3123, N3121, N3071);
or OR2 (N3124, N3116, N694);
xor XOR2 (N3125, N3114, N2681);
xor XOR2 (N3126, N3106, N857);
not NOT1 (N3127, N3117);
or OR2 (N3128, N3127, N2965);
and AND3 (N3129, N3113, N2230, N1814);
nand NAND2 (N3130, N3128, N1132);
buf BUF1 (N3131, N3126);
nor NOR4 (N3132, N3118, N1035, N1492, N244);
buf BUF1 (N3133, N3131);
nand NAND2 (N3134, N3133, N2116);
not NOT1 (N3135, N3122);
buf BUF1 (N3136, N3135);
and AND4 (N3137, N3124, N2172, N1901, N2002);
and AND2 (N3138, N3125, N728);
nor NOR2 (N3139, N3138, N407);
not NOT1 (N3140, N3132);
xor XOR2 (N3141, N3123, N252);
nor NOR3 (N3142, N3090, N173, N320);
nand NAND3 (N3143, N3130, N1013, N2705);
buf BUF1 (N3144, N3143);
nor NOR3 (N3145, N3119, N3101, N2619);
not NOT1 (N3146, N3129);
and AND4 (N3147, N3142, N2899, N862, N1665);
not NOT1 (N3148, N3144);
or OR2 (N3149, N3148, N1570);
buf BUF1 (N3150, N3134);
nand NAND4 (N3151, N3147, N2217, N1124, N1419);
and AND3 (N3152, N3140, N25, N1841);
not NOT1 (N3153, N3139);
not NOT1 (N3154, N3150);
buf BUF1 (N3155, N3152);
or OR3 (N3156, N3136, N805, N3091);
xor XOR2 (N3157, N3153, N1671);
and AND3 (N3158, N3145, N2134, N2544);
or OR2 (N3159, N3137, N1400);
xor XOR2 (N3160, N3158, N2035);
nor NOR3 (N3161, N3146, N2648, N631);
nand NAND3 (N3162, N3141, N3050, N2005);
and AND2 (N3163, N3149, N2624);
xor XOR2 (N3164, N3162, N2397);
not NOT1 (N3165, N3164);
not NOT1 (N3166, N3151);
nand NAND4 (N3167, N3160, N2919, N1511, N390);
xor XOR2 (N3168, N3159, N1952);
buf BUF1 (N3169, N3155);
or OR3 (N3170, N3165, N2585, N2381);
xor XOR2 (N3171, N3157, N1342);
xor XOR2 (N3172, N3169, N1473);
buf BUF1 (N3173, N3156);
and AND3 (N3174, N3161, N1066, N1720);
xor XOR2 (N3175, N3172, N2185);
nor NOR2 (N3176, N3175, N2226);
or OR3 (N3177, N3166, N105, N2360);
buf BUF1 (N3178, N3177);
nand NAND2 (N3179, N3167, N2389);
buf BUF1 (N3180, N3168);
nor NOR4 (N3181, N3179, N3037, N1892, N1474);
xor XOR2 (N3182, N3178, N1594);
and AND3 (N3183, N3171, N3086, N2364);
or OR4 (N3184, N3180, N1243, N3035, N3155);
and AND4 (N3185, N3184, N690, N1903, N920);
not NOT1 (N3186, N3181);
or OR3 (N3187, N3170, N642, N890);
xor XOR2 (N3188, N3186, N658);
and AND3 (N3189, N3185, N3160, N108);
nand NAND3 (N3190, N3163, N1005, N1900);
nand NAND2 (N3191, N3174, N161);
nor NOR2 (N3192, N3154, N1545);
nor NOR3 (N3193, N3191, N1821, N1265);
xor XOR2 (N3194, N3188, N2531);
nor NOR2 (N3195, N3187, N2069);
or OR2 (N3196, N3183, N2900);
nand NAND2 (N3197, N3195, N2984);
and AND3 (N3198, N3193, N1058, N2232);
not NOT1 (N3199, N3189);
not NOT1 (N3200, N3197);
xor XOR2 (N3201, N3194, N410);
nand NAND2 (N3202, N3200, N3054);
nor NOR4 (N3203, N3192, N2156, N1468, N931);
nor NOR4 (N3204, N3176, N1519, N1571, N1210);
nand NAND3 (N3205, N3201, N482, N1985);
not NOT1 (N3206, N3205);
buf BUF1 (N3207, N3198);
xor XOR2 (N3208, N3190, N2174);
or OR4 (N3209, N3204, N12, N1623, N1363);
buf BUF1 (N3210, N3182);
nand NAND3 (N3211, N3196, N808, N3208);
or OR4 (N3212, N1410, N1819, N2547, N2587);
or OR2 (N3213, N3211, N76);
and AND3 (N3214, N3210, N991, N2738);
buf BUF1 (N3215, N3207);
nand NAND4 (N3216, N3212, N1023, N1991, N33);
or OR3 (N3217, N3206, N699, N711);
nor NOR2 (N3218, N3202, N2232);
buf BUF1 (N3219, N3203);
not NOT1 (N3220, N3216);
buf BUF1 (N3221, N3173);
not NOT1 (N3222, N3215);
nor NOR4 (N3223, N3218, N3055, N2965, N111);
not NOT1 (N3224, N3221);
not NOT1 (N3225, N3219);
not NOT1 (N3226, N3209);
nor NOR2 (N3227, N3222, N3023);
nand NAND4 (N3228, N3227, N230, N3049, N1096);
or OR4 (N3229, N3224, N1209, N1873, N607);
and AND4 (N3230, N3213, N384, N783, N1988);
and AND2 (N3231, N3223, N121);
not NOT1 (N3232, N3199);
buf BUF1 (N3233, N3226);
and AND4 (N3234, N3229, N1154, N3070, N2142);
not NOT1 (N3235, N3234);
nor NOR3 (N3236, N3214, N1010, N1884);
and AND4 (N3237, N3217, N10, N1761, N2996);
or OR4 (N3238, N3233, N2710, N1936, N2561);
nand NAND4 (N3239, N3237, N71, N1335, N97);
or OR2 (N3240, N3228, N565);
buf BUF1 (N3241, N3236);
nand NAND4 (N3242, N3240, N515, N745, N2349);
and AND4 (N3243, N3220, N2435, N2360, N1570);
buf BUF1 (N3244, N3241);
or OR3 (N3245, N3231, N755, N2412);
and AND2 (N3246, N3225, N2720);
not NOT1 (N3247, N3239);
nor NOR2 (N3248, N3238, N2235);
or OR3 (N3249, N3246, N3229, N1406);
nor NOR3 (N3250, N3242, N2611, N1984);
nand NAND4 (N3251, N3249, N1158, N1688, N826);
not NOT1 (N3252, N3250);
xor XOR2 (N3253, N3230, N1603);
buf BUF1 (N3254, N3248);
or OR3 (N3255, N3247, N2369, N613);
and AND2 (N3256, N3232, N2201);
xor XOR2 (N3257, N3252, N1720);
nor NOR3 (N3258, N3255, N2439, N581);
nand NAND4 (N3259, N3253, N1203, N2226, N516);
xor XOR2 (N3260, N3258, N984);
not NOT1 (N3261, N3254);
nor NOR2 (N3262, N3245, N1943);
or OR2 (N3263, N3260, N2796);
and AND3 (N3264, N3235, N1956, N215);
nand NAND3 (N3265, N3263, N2263, N347);
not NOT1 (N3266, N3243);
and AND4 (N3267, N3264, N1155, N1929, N594);
not NOT1 (N3268, N3261);
nand NAND4 (N3269, N3251, N2220, N1503, N1052);
and AND4 (N3270, N3267, N2542, N2811, N1397);
and AND2 (N3271, N3259, N302);
nor NOR3 (N3272, N3257, N1603, N1825);
buf BUF1 (N3273, N3266);
buf BUF1 (N3274, N3271);
nand NAND2 (N3275, N3256, N534);
nor NOR2 (N3276, N3268, N2749);
or OR4 (N3277, N3273, N1275, N1128, N2603);
xor XOR2 (N3278, N3276, N881);
nand NAND2 (N3279, N3274, N205);
not NOT1 (N3280, N3279);
not NOT1 (N3281, N3262);
buf BUF1 (N3282, N3269);
nor NOR2 (N3283, N3270, N3084);
and AND3 (N3284, N3277, N3215, N2340);
nor NOR4 (N3285, N3284, N2603, N2025, N2433);
and AND2 (N3286, N3265, N1326);
buf BUF1 (N3287, N3272);
or OR4 (N3288, N3282, N1840, N374, N882);
nand NAND4 (N3289, N3280, N2956, N40, N327);
not NOT1 (N3290, N3275);
buf BUF1 (N3291, N3288);
or OR2 (N3292, N3289, N3148);
nor NOR4 (N3293, N3281, N1420, N739, N2065);
nand NAND2 (N3294, N3292, N1035);
xor XOR2 (N3295, N3290, N148);
buf BUF1 (N3296, N3293);
and AND4 (N3297, N3278, N1004, N1714, N3275);
and AND2 (N3298, N3297, N2916);
not NOT1 (N3299, N3287);
and AND2 (N3300, N3299, N2691);
or OR3 (N3301, N3298, N1254, N536);
nand NAND4 (N3302, N3286, N1845, N48, N2805);
or OR3 (N3303, N3291, N2528, N2379);
not NOT1 (N3304, N3285);
or OR2 (N3305, N3303, N1487);
nor NOR3 (N3306, N3301, N2519, N3062);
xor XOR2 (N3307, N3283, N3221);
and AND3 (N3308, N3307, N1417, N2601);
xor XOR2 (N3309, N3244, N2286);
or OR2 (N3310, N3304, N2799);
not NOT1 (N3311, N3294);
xor XOR2 (N3312, N3296, N1307);
nor NOR4 (N3313, N3312, N325, N358, N2851);
nor NOR3 (N3314, N3300, N1985, N2286);
nor NOR3 (N3315, N3309, N230, N665);
and AND3 (N3316, N3305, N2995, N1331);
nor NOR2 (N3317, N3313, N1780);
nor NOR4 (N3318, N3314, N1977, N2100, N2085);
and AND4 (N3319, N3317, N2620, N2071, N286);
buf BUF1 (N3320, N3315);
not NOT1 (N3321, N3320);
xor XOR2 (N3322, N3308, N2091);
xor XOR2 (N3323, N3311, N861);
and AND3 (N3324, N3318, N1619, N205);
and AND4 (N3325, N3316, N2523, N2014, N2704);
and AND3 (N3326, N3306, N744, N2516);
buf BUF1 (N3327, N3319);
xor XOR2 (N3328, N3324, N1261);
nand NAND2 (N3329, N3323, N2337);
nand NAND2 (N3330, N3325, N2508);
or OR4 (N3331, N3302, N2964, N3272, N917);
buf BUF1 (N3332, N3327);
xor XOR2 (N3333, N3328, N1122);
nor NOR2 (N3334, N3333, N1695);
and AND4 (N3335, N3330, N1982, N3092, N272);
xor XOR2 (N3336, N3295, N2272);
nor NOR3 (N3337, N3336, N3154, N136);
and AND4 (N3338, N3334, N2832, N1604, N1744);
not NOT1 (N3339, N3337);
not NOT1 (N3340, N3332);
and AND3 (N3341, N3340, N835, N2796);
and AND4 (N3342, N3331, N368, N895, N2032);
buf BUF1 (N3343, N3321);
or OR3 (N3344, N3329, N982, N2627);
nand NAND3 (N3345, N3344, N2013, N3318);
xor XOR2 (N3346, N3345, N2376);
and AND2 (N3347, N3335, N832);
and AND4 (N3348, N3346, N2456, N3038, N207);
buf BUF1 (N3349, N3338);
not NOT1 (N3350, N3342);
nor NOR2 (N3351, N3350, N983);
buf BUF1 (N3352, N3339);
or OR4 (N3353, N3349, N708, N2147, N2585);
xor XOR2 (N3354, N3341, N3208);
or OR2 (N3355, N3354, N2457);
not NOT1 (N3356, N3353);
not NOT1 (N3357, N3356);
nand NAND4 (N3358, N3347, N359, N1802, N1325);
and AND4 (N3359, N3352, N838, N2126, N911);
nand NAND2 (N3360, N3357, N694);
not NOT1 (N3361, N3360);
and AND3 (N3362, N3358, N1481, N186);
nand NAND3 (N3363, N3362, N1311, N1855);
and AND4 (N3364, N3351, N3111, N1384, N2570);
nor NOR2 (N3365, N3326, N352);
buf BUF1 (N3366, N3365);
xor XOR2 (N3367, N3364, N2283);
xor XOR2 (N3368, N3367, N3153);
nor NOR3 (N3369, N3359, N3168, N1774);
or OR3 (N3370, N3322, N383, N1107);
buf BUF1 (N3371, N3361);
xor XOR2 (N3372, N3363, N107);
xor XOR2 (N3373, N3343, N1887);
not NOT1 (N3374, N3370);
and AND2 (N3375, N3368, N3362);
buf BUF1 (N3376, N3310);
nor NOR3 (N3377, N3376, N2671, N3168);
not NOT1 (N3378, N3348);
nand NAND3 (N3379, N3375, N2751, N3331);
nor NOR4 (N3380, N3374, N1321, N512, N413);
or OR2 (N3381, N3380, N1686);
nand NAND4 (N3382, N3366, N3029, N2064, N2968);
buf BUF1 (N3383, N3373);
nand NAND4 (N3384, N3379, N2493, N3199, N1541);
nor NOR4 (N3385, N3355, N628, N2972, N1208);
xor XOR2 (N3386, N3384, N62);
and AND4 (N3387, N3377, N2015, N2215, N3348);
nand NAND2 (N3388, N3386, N1219);
xor XOR2 (N3389, N3385, N2856);
nand NAND2 (N3390, N3389, N1481);
and AND3 (N3391, N3387, N2732, N2702);
buf BUF1 (N3392, N3371);
and AND2 (N3393, N3388, N519);
nand NAND3 (N3394, N3391, N1701, N1656);
nand NAND4 (N3395, N3372, N1458, N2865, N622);
nor NOR4 (N3396, N3392, N429, N645, N700);
nor NOR2 (N3397, N3383, N256);
and AND3 (N3398, N3393, N2313, N2584);
nand NAND3 (N3399, N3378, N2038, N1561);
and AND2 (N3400, N3399, N2663);
nor NOR3 (N3401, N3398, N1102, N3116);
not NOT1 (N3402, N3369);
or OR2 (N3403, N3400, N214);
nand NAND2 (N3404, N3381, N3279);
nor NOR4 (N3405, N3404, N2042, N717, N1689);
nand NAND2 (N3406, N3394, N2917);
not NOT1 (N3407, N3402);
not NOT1 (N3408, N3382);
not NOT1 (N3409, N3406);
nor NOR4 (N3410, N3408, N3323, N2301, N2346);
nand NAND2 (N3411, N3395, N3281);
and AND3 (N3412, N3396, N2666, N2994);
xor XOR2 (N3413, N3411, N2072);
and AND2 (N3414, N3409, N2349);
nor NOR4 (N3415, N3410, N1299, N1225, N3131);
or OR3 (N3416, N3390, N3080, N2953);
xor XOR2 (N3417, N3412, N1877);
and AND4 (N3418, N3414, N516, N367, N1362);
and AND3 (N3419, N3397, N2310, N1469);
nand NAND2 (N3420, N3417, N477);
buf BUF1 (N3421, N3420);
xor XOR2 (N3422, N3419, N2202);
nor NOR3 (N3423, N3405, N2082, N2962);
nand NAND2 (N3424, N3423, N3038);
nand NAND4 (N3425, N3401, N2183, N2610, N1843);
or OR2 (N3426, N3413, N985);
and AND4 (N3427, N3421, N680, N860, N3420);
xor XOR2 (N3428, N3416, N2071);
buf BUF1 (N3429, N3403);
nor NOR2 (N3430, N3424, N1980);
nor NOR2 (N3431, N3426, N162);
xor XOR2 (N3432, N3425, N2468);
and AND3 (N3433, N3427, N579, N804);
buf BUF1 (N3434, N3431);
xor XOR2 (N3435, N3418, N1658);
and AND3 (N3436, N3407, N286, N723);
nor NOR3 (N3437, N3435, N3166, N957);
xor XOR2 (N3438, N3415, N1545);
or OR4 (N3439, N3430, N2318, N223, N2510);
xor XOR2 (N3440, N3438, N1792);
or OR2 (N3441, N3434, N514);
nand NAND4 (N3442, N3437, N2644, N1381, N3033);
xor XOR2 (N3443, N3442, N2915);
xor XOR2 (N3444, N3439, N388);
and AND3 (N3445, N3433, N1419, N1434);
nand NAND4 (N3446, N3445, N1970, N271, N1539);
nor NOR2 (N3447, N3436, N2461);
buf BUF1 (N3448, N3440);
and AND3 (N3449, N3443, N258, N1894);
not NOT1 (N3450, N3444);
or OR2 (N3451, N3448, N2414);
xor XOR2 (N3452, N3422, N1860);
nor NOR4 (N3453, N3432, N1695, N1336, N3214);
nor NOR3 (N3454, N3450, N3405, N2629);
nand NAND4 (N3455, N3449, N2836, N1639, N1933);
nand NAND4 (N3456, N3446, N2147, N3073, N1720);
buf BUF1 (N3457, N3441);
and AND3 (N3458, N3456, N2703, N1669);
and AND2 (N3459, N3452, N515);
and AND4 (N3460, N3447, N131, N1172, N3036);
xor XOR2 (N3461, N3453, N1832);
buf BUF1 (N3462, N3454);
and AND4 (N3463, N3455, N789, N2375, N2004);
nor NOR2 (N3464, N3461, N3107);
or OR2 (N3465, N3464, N2608);
xor XOR2 (N3466, N3429, N2425);
xor XOR2 (N3467, N3462, N2306);
xor XOR2 (N3468, N3428, N1092);
xor XOR2 (N3469, N3466, N371);
not NOT1 (N3470, N3468);
or OR3 (N3471, N3459, N633, N1137);
buf BUF1 (N3472, N3451);
buf BUF1 (N3473, N3457);
and AND3 (N3474, N3460, N3349, N2828);
not NOT1 (N3475, N3474);
not NOT1 (N3476, N3475);
and AND3 (N3477, N3471, N1592, N3110);
buf BUF1 (N3478, N3476);
buf BUF1 (N3479, N3477);
and AND4 (N3480, N3458, N933, N3430, N2076);
not NOT1 (N3481, N3472);
not NOT1 (N3482, N3480);
nor NOR4 (N3483, N3463, N3326, N2550, N3007);
nor NOR4 (N3484, N3473, N2977, N2640, N990);
or OR4 (N3485, N3481, N2322, N918, N3407);
and AND3 (N3486, N3465, N1931, N2107);
or OR2 (N3487, N3486, N834);
and AND4 (N3488, N3478, N1699, N2818, N2334);
or OR4 (N3489, N3485, N1935, N1033, N26);
or OR4 (N3490, N3470, N3088, N3329, N2282);
buf BUF1 (N3491, N3489);
and AND2 (N3492, N3488, N2293);
or OR2 (N3493, N3483, N1175);
nor NOR3 (N3494, N3469, N2624, N2814);
xor XOR2 (N3495, N3491, N1410);
and AND4 (N3496, N3482, N2532, N2735, N1719);
and AND3 (N3497, N3487, N2758, N2945);
nor NOR4 (N3498, N3495, N492, N3117, N1562);
xor XOR2 (N3499, N3467, N1162);
nand NAND2 (N3500, N3494, N1479);
buf BUF1 (N3501, N3479);
nor NOR4 (N3502, N3496, N1368, N1806, N48);
nor NOR3 (N3503, N3501, N3046, N3028);
xor XOR2 (N3504, N3500, N1820);
not NOT1 (N3505, N3504);
or OR2 (N3506, N3492, N961);
nand NAND3 (N3507, N3506, N1057, N1663);
buf BUF1 (N3508, N3505);
xor XOR2 (N3509, N3484, N1092);
not NOT1 (N3510, N3503);
buf BUF1 (N3511, N3499);
nor NOR4 (N3512, N3507, N766, N768, N1387);
or OR2 (N3513, N3490, N2);
buf BUF1 (N3514, N3498);
and AND2 (N3515, N3513, N1905);
buf BUF1 (N3516, N3510);
or OR3 (N3517, N3516, N3382, N2840);
buf BUF1 (N3518, N3509);
or OR3 (N3519, N3497, N1581, N1619);
not NOT1 (N3520, N3519);
and AND2 (N3521, N3515, N117);
or OR4 (N3522, N3517, N743, N2476, N437);
not NOT1 (N3523, N3514);
xor XOR2 (N3524, N3502, N1345);
or OR4 (N3525, N3493, N173, N1993, N3389);
or OR2 (N3526, N3521, N592);
buf BUF1 (N3527, N3524);
xor XOR2 (N3528, N3512, N595);
not NOT1 (N3529, N3518);
buf BUF1 (N3530, N3522);
buf BUF1 (N3531, N3511);
not NOT1 (N3532, N3528);
nand NAND2 (N3533, N3531, N1553);
and AND3 (N3534, N3532, N8, N2913);
not NOT1 (N3535, N3520);
buf BUF1 (N3536, N3526);
not NOT1 (N3537, N3523);
or OR2 (N3538, N3529, N479);
not NOT1 (N3539, N3530);
and AND2 (N3540, N3533, N1757);
buf BUF1 (N3541, N3538);
buf BUF1 (N3542, N3540);
nand NAND4 (N3543, N3537, N1646, N2341, N2383);
nor NOR3 (N3544, N3539, N2882, N2319);
buf BUF1 (N3545, N3536);
buf BUF1 (N3546, N3527);
not NOT1 (N3547, N3545);
buf BUF1 (N3548, N3534);
or OR2 (N3549, N3525, N2106);
and AND2 (N3550, N3535, N2275);
not NOT1 (N3551, N3547);
not NOT1 (N3552, N3551);
buf BUF1 (N3553, N3550);
buf BUF1 (N3554, N3549);
nor NOR4 (N3555, N3544, N3414, N1080, N2448);
and AND3 (N3556, N3548, N1111, N3041);
nor NOR2 (N3557, N3543, N2245);
not NOT1 (N3558, N3542);
and AND3 (N3559, N3546, N884, N268);
not NOT1 (N3560, N3556);
nand NAND3 (N3561, N3508, N834, N2931);
nor NOR4 (N3562, N3552, N2922, N425, N3327);
xor XOR2 (N3563, N3557, N943);
nor NOR2 (N3564, N3555, N307);
and AND4 (N3565, N3541, N1303, N3455, N79);
nand NAND2 (N3566, N3565, N789);
buf BUF1 (N3567, N3561);
xor XOR2 (N3568, N3567, N3265);
buf BUF1 (N3569, N3558);
buf BUF1 (N3570, N3566);
buf BUF1 (N3571, N3570);
or OR3 (N3572, N3563, N2383, N2542);
or OR4 (N3573, N3569, N1595, N2267, N1580);
not NOT1 (N3574, N3568);
xor XOR2 (N3575, N3560, N3500);
not NOT1 (N3576, N3574);
not NOT1 (N3577, N3564);
buf BUF1 (N3578, N3575);
or OR2 (N3579, N3573, N1114);
buf BUF1 (N3580, N3579);
nor NOR4 (N3581, N3580, N1716, N592, N3465);
not NOT1 (N3582, N3576);
not NOT1 (N3583, N3578);
nand NAND4 (N3584, N3554, N2928, N3182, N987);
buf BUF1 (N3585, N3577);
buf BUF1 (N3586, N3562);
nand NAND3 (N3587, N3584, N1737, N2871);
not NOT1 (N3588, N3586);
and AND4 (N3589, N3572, N1096, N2927, N186);
nor NOR4 (N3590, N3589, N2639, N142, N1649);
nor NOR4 (N3591, N3571, N2995, N1066, N553);
nand NAND2 (N3592, N3581, N972);
buf BUF1 (N3593, N3553);
buf BUF1 (N3594, N3593);
and AND4 (N3595, N3559, N3160, N2120, N1313);
not NOT1 (N3596, N3595);
nor NOR4 (N3597, N3594, N1087, N2313, N701);
nand NAND3 (N3598, N3591, N1558, N1165);
not NOT1 (N3599, N3596);
or OR2 (N3600, N3598, N2277);
not NOT1 (N3601, N3590);
and AND4 (N3602, N3582, N2064, N3572, N430);
nor NOR3 (N3603, N3587, N424, N1574);
xor XOR2 (N3604, N3597, N1839);
nand NAND2 (N3605, N3603, N320);
xor XOR2 (N3606, N3600, N2410);
nand NAND4 (N3607, N3592, N2291, N471, N1614);
nor NOR4 (N3608, N3607, N2565, N685, N1193);
xor XOR2 (N3609, N3602, N533);
not NOT1 (N3610, N3605);
and AND3 (N3611, N3585, N3166, N2584);
nor NOR4 (N3612, N3604, N2748, N3305, N3463);
buf BUF1 (N3613, N3599);
nand NAND2 (N3614, N3610, N2942);
or OR2 (N3615, N3613, N437);
or OR2 (N3616, N3615, N996);
nor NOR4 (N3617, N3601, N286, N3571, N2918);
nand NAND4 (N3618, N3588, N796, N2564, N918);
xor XOR2 (N3619, N3609, N2339);
nand NAND3 (N3620, N3608, N2354, N2085);
not NOT1 (N3621, N3620);
or OR3 (N3622, N3614, N2671, N2694);
buf BUF1 (N3623, N3621);
buf BUF1 (N3624, N3616);
or OR3 (N3625, N3618, N2608, N2155);
xor XOR2 (N3626, N3611, N80);
and AND3 (N3627, N3617, N979, N1065);
or OR2 (N3628, N3625, N1266);
xor XOR2 (N3629, N3583, N2776);
xor XOR2 (N3630, N3606, N2065);
xor XOR2 (N3631, N3619, N3334);
nor NOR3 (N3632, N3612, N1340, N2428);
not NOT1 (N3633, N3630);
nand NAND3 (N3634, N3624, N3348, N2294);
nor NOR2 (N3635, N3629, N1803);
xor XOR2 (N3636, N3628, N850);
or OR4 (N3637, N3627, N402, N1479, N1689);
nor NOR3 (N3638, N3637, N2322, N3421);
nand NAND4 (N3639, N3623, N529, N3062, N1306);
or OR4 (N3640, N3632, N968, N1006, N2479);
not NOT1 (N3641, N3640);
and AND2 (N3642, N3635, N2678);
nand NAND4 (N3643, N3636, N2591, N2302, N2749);
buf BUF1 (N3644, N3643);
and AND2 (N3645, N3638, N1811);
buf BUF1 (N3646, N3642);
not NOT1 (N3647, N3631);
or OR4 (N3648, N3641, N1895, N2086, N549);
nor NOR3 (N3649, N3622, N2422, N2380);
xor XOR2 (N3650, N3648, N2498);
and AND2 (N3651, N3646, N424);
nand NAND4 (N3652, N3645, N2481, N1013, N3473);
buf BUF1 (N3653, N3651);
not NOT1 (N3654, N3647);
or OR4 (N3655, N3633, N450, N2609, N2504);
and AND4 (N3656, N3654, N1688, N2617, N2087);
xor XOR2 (N3657, N3639, N1543);
and AND3 (N3658, N3626, N979, N1910);
buf BUF1 (N3659, N3644);
xor XOR2 (N3660, N3650, N110);
nor NOR3 (N3661, N3656, N475, N2365);
nand NAND2 (N3662, N3659, N3388);
and AND4 (N3663, N3649, N208, N1217, N3174);
nand NAND2 (N3664, N3653, N3286);
nand NAND4 (N3665, N3662, N1945, N930, N1784);
and AND4 (N3666, N3665, N2290, N1706, N480);
nor NOR3 (N3667, N3652, N2327, N2949);
buf BUF1 (N3668, N3634);
xor XOR2 (N3669, N3664, N1986);
buf BUF1 (N3670, N3666);
nand NAND4 (N3671, N3667, N1951, N550, N353);
and AND2 (N3672, N3663, N1310);
nor NOR4 (N3673, N3660, N529, N2036, N3383);
or OR3 (N3674, N3668, N478, N927);
nor NOR4 (N3675, N3671, N2374, N3111, N3031);
xor XOR2 (N3676, N3655, N3576);
and AND3 (N3677, N3674, N93, N3169);
and AND2 (N3678, N3676, N2372);
and AND3 (N3679, N3677, N3677, N2514);
nand NAND3 (N3680, N3658, N1498, N2918);
and AND4 (N3681, N3657, N2170, N155, N926);
nor NOR2 (N3682, N3669, N37);
or OR4 (N3683, N3672, N1143, N2080, N2812);
xor XOR2 (N3684, N3681, N2281);
buf BUF1 (N3685, N3680);
nand NAND2 (N3686, N3673, N1163);
nor NOR3 (N3687, N3683, N2590, N3136);
nand NAND2 (N3688, N3682, N885);
buf BUF1 (N3689, N3688);
or OR3 (N3690, N3684, N782, N401);
nand NAND4 (N3691, N3689, N2702, N1137, N957);
buf BUF1 (N3692, N3679);
and AND2 (N3693, N3675, N1741);
xor XOR2 (N3694, N3690, N3027);
xor XOR2 (N3695, N3678, N597);
nor NOR4 (N3696, N3695, N2596, N1934, N2610);
or OR2 (N3697, N3685, N1475);
nor NOR3 (N3698, N3692, N2708, N3295);
or OR2 (N3699, N3694, N3302);
and AND3 (N3700, N3699, N645, N343);
nor NOR2 (N3701, N3693, N1070);
nand NAND3 (N3702, N3661, N2836, N1798);
nor NOR4 (N3703, N3701, N121, N787, N2145);
and AND3 (N3704, N3702, N2881, N3377);
not NOT1 (N3705, N3686);
buf BUF1 (N3706, N3698);
or OR2 (N3707, N3697, N765);
not NOT1 (N3708, N3696);
or OR4 (N3709, N3687, N2255, N2825, N2544);
nand NAND2 (N3710, N3700, N2555);
or OR2 (N3711, N3707, N2742);
xor XOR2 (N3712, N3710, N3184);
xor XOR2 (N3713, N3703, N3673);
or OR4 (N3714, N3706, N3521, N2296, N1734);
or OR3 (N3715, N3670, N2728, N2317);
buf BUF1 (N3716, N3711);
buf BUF1 (N3717, N3704);
nor NOR4 (N3718, N3705, N126, N807, N1725);
buf BUF1 (N3719, N3712);
buf BUF1 (N3720, N3713);
nand NAND4 (N3721, N3709, N864, N957, N3687);
or OR2 (N3722, N3721, N933);
buf BUF1 (N3723, N3719);
and AND3 (N3724, N3691, N3631, N2640);
buf BUF1 (N3725, N3723);
not NOT1 (N3726, N3718);
buf BUF1 (N3727, N3708);
buf BUF1 (N3728, N3724);
buf BUF1 (N3729, N3716);
or OR2 (N3730, N3729, N1624);
buf BUF1 (N3731, N3717);
nor NOR4 (N3732, N3714, N3660, N2319, N3037);
and AND2 (N3733, N3731, N3600);
and AND3 (N3734, N3733, N203, N2733);
or OR3 (N3735, N3720, N2179, N2173);
and AND3 (N3736, N3722, N524, N2007);
and AND3 (N3737, N3734, N81, N2167);
nand NAND3 (N3738, N3727, N2737, N1176);
nor NOR4 (N3739, N3737, N1725, N2198, N3731);
buf BUF1 (N3740, N3732);
buf BUF1 (N3741, N3726);
and AND3 (N3742, N3730, N1804, N127);
and AND2 (N3743, N3739, N1950);
nand NAND2 (N3744, N3740, N3590);
not NOT1 (N3745, N3715);
nand NAND4 (N3746, N3744, N3258, N892, N2852);
buf BUF1 (N3747, N3745);
and AND4 (N3748, N3735, N2295, N3435, N2419);
and AND2 (N3749, N3742, N2145);
nand NAND2 (N3750, N3747, N2148);
nor NOR4 (N3751, N3748, N3646, N3209, N709);
and AND2 (N3752, N3750, N1905);
xor XOR2 (N3753, N3736, N3035);
nand NAND2 (N3754, N3743, N930);
not NOT1 (N3755, N3753);
xor XOR2 (N3756, N3728, N1999);
or OR2 (N3757, N3741, N481);
or OR2 (N3758, N3725, N3315);
nor NOR2 (N3759, N3746, N3321);
xor XOR2 (N3760, N3756, N241);
nor NOR2 (N3761, N3749, N2917);
xor XOR2 (N3762, N3738, N1556);
or OR4 (N3763, N3755, N301, N691, N562);
and AND3 (N3764, N3763, N2663, N2903);
and AND2 (N3765, N3760, N1141);
and AND2 (N3766, N3752, N3734);
not NOT1 (N3767, N3762);
nor NOR2 (N3768, N3758, N833);
buf BUF1 (N3769, N3759);
xor XOR2 (N3770, N3765, N209);
buf BUF1 (N3771, N3751);
nand NAND4 (N3772, N3757, N1026, N2339, N3423);
or OR3 (N3773, N3770, N119, N241);
and AND4 (N3774, N3769, N2700, N1436, N737);
or OR4 (N3775, N3768, N3542, N903, N2986);
not NOT1 (N3776, N3772);
and AND3 (N3777, N3766, N2271, N3695);
not NOT1 (N3778, N3761);
nand NAND2 (N3779, N3776, N616);
not NOT1 (N3780, N3767);
nand NAND3 (N3781, N3764, N734, N2109);
and AND2 (N3782, N3771, N1108);
buf BUF1 (N3783, N3773);
nor NOR4 (N3784, N3782, N3753, N272, N3456);
buf BUF1 (N3785, N3780);
nand NAND3 (N3786, N3774, N405, N3);
nor NOR3 (N3787, N3783, N2338, N1913);
and AND4 (N3788, N3786, N1051, N2573, N3533);
buf BUF1 (N3789, N3787);
or OR2 (N3790, N3789, N2661);
nand NAND4 (N3791, N3777, N3011, N2261, N2990);
not NOT1 (N3792, N3784);
or OR3 (N3793, N3790, N1432, N1590);
buf BUF1 (N3794, N3793);
nand NAND3 (N3795, N3775, N2880, N1067);
buf BUF1 (N3796, N3754);
and AND3 (N3797, N3792, N149, N2161);
nand NAND3 (N3798, N3795, N1631, N1780);
and AND2 (N3799, N3796, N1661);
and AND4 (N3800, N3778, N2902, N951, N3288);
buf BUF1 (N3801, N3781);
xor XOR2 (N3802, N3791, N2648);
nor NOR2 (N3803, N3779, N3213);
buf BUF1 (N3804, N3803);
nand NAND3 (N3805, N3785, N943, N3519);
xor XOR2 (N3806, N3800, N1372);
nand NAND3 (N3807, N3788, N2819, N2227);
or OR2 (N3808, N3802, N3800);
nor NOR4 (N3809, N3797, N1302, N350, N3232);
and AND2 (N3810, N3804, N613);
nand NAND2 (N3811, N3799, N40);
and AND2 (N3812, N3798, N903);
not NOT1 (N3813, N3805);
xor XOR2 (N3814, N3801, N193);
or OR3 (N3815, N3808, N49, N3705);
or OR4 (N3816, N3814, N1521, N3783, N3439);
buf BUF1 (N3817, N3815);
and AND3 (N3818, N3816, N3297, N1457);
buf BUF1 (N3819, N3817);
xor XOR2 (N3820, N3818, N2611);
nor NOR4 (N3821, N3819, N3796, N861, N2423);
xor XOR2 (N3822, N3811, N1409);
or OR2 (N3823, N3810, N885);
nor NOR3 (N3824, N3821, N1573, N928);
not NOT1 (N3825, N3794);
buf BUF1 (N3826, N3822);
nor NOR4 (N3827, N3825, N2449, N2304, N123);
xor XOR2 (N3828, N3827, N1255);
buf BUF1 (N3829, N3806);
xor XOR2 (N3830, N3807, N604);
not NOT1 (N3831, N3813);
or OR4 (N3832, N3824, N3427, N1682, N3306);
buf BUF1 (N3833, N3820);
or OR3 (N3834, N3829, N3155, N1411);
xor XOR2 (N3835, N3831, N1284);
or OR3 (N3836, N3835, N1205, N27);
or OR3 (N3837, N3828, N1413, N204);
nor NOR3 (N3838, N3809, N2476, N2104);
nor NOR4 (N3839, N3838, N2853, N2859, N1893);
and AND3 (N3840, N3812, N2068, N3158);
or OR2 (N3841, N3830, N882);
xor XOR2 (N3842, N3840, N3147);
nor NOR2 (N3843, N3834, N1076);
nor NOR3 (N3844, N3841, N2859, N2078);
and AND2 (N3845, N3832, N3656);
buf BUF1 (N3846, N3839);
nand NAND3 (N3847, N3844, N535, N755);
not NOT1 (N3848, N3833);
and AND4 (N3849, N3837, N1117, N1570, N760);
buf BUF1 (N3850, N3836);
nor NOR4 (N3851, N3849, N1001, N1001, N3593);
nand NAND2 (N3852, N3846, N610);
nand NAND4 (N3853, N3852, N931, N2196, N2363);
and AND2 (N3854, N3853, N1755);
or OR3 (N3855, N3845, N3603, N731);
not NOT1 (N3856, N3851);
buf BUF1 (N3857, N3856);
or OR3 (N3858, N3857, N498, N983);
xor XOR2 (N3859, N3858, N2025);
nand NAND2 (N3860, N3855, N2186);
nand NAND3 (N3861, N3860, N583, N1573);
not NOT1 (N3862, N3842);
and AND2 (N3863, N3850, N1506);
or OR4 (N3864, N3823, N3457, N3078, N2664);
nand NAND4 (N3865, N3848, N3444, N1392, N807);
not NOT1 (N3866, N3826);
or OR2 (N3867, N3864, N2616);
nand NAND4 (N3868, N3859, N1261, N3161, N2503);
nand NAND4 (N3869, N3847, N2407, N259, N16);
nor NOR2 (N3870, N3865, N322);
buf BUF1 (N3871, N3869);
or OR3 (N3872, N3868, N1194, N3770);
not NOT1 (N3873, N3862);
buf BUF1 (N3874, N3863);
xor XOR2 (N3875, N3871, N257);
xor XOR2 (N3876, N3874, N2446);
xor XOR2 (N3877, N3866, N3380);
buf BUF1 (N3878, N3870);
xor XOR2 (N3879, N3873, N2342);
and AND4 (N3880, N3878, N3142, N119, N2083);
nor NOR3 (N3881, N3880, N1127, N1778);
or OR3 (N3882, N3867, N1570, N1482);
or OR2 (N3883, N3881, N3528);
and AND4 (N3884, N3843, N3506, N1491, N1826);
and AND2 (N3885, N3882, N3398);
nand NAND4 (N3886, N3854, N1381, N1652, N1834);
and AND2 (N3887, N3876, N616);
and AND4 (N3888, N3887, N2223, N606, N1607);
xor XOR2 (N3889, N3877, N2753);
nor NOR2 (N3890, N3872, N1700);
not NOT1 (N3891, N3879);
nor NOR4 (N3892, N3875, N560, N2008, N567);
not NOT1 (N3893, N3891);
and AND4 (N3894, N3886, N1276, N956, N750);
xor XOR2 (N3895, N3893, N3557);
nor NOR3 (N3896, N3895, N3808, N2843);
not NOT1 (N3897, N3883);
and AND2 (N3898, N3889, N3872);
not NOT1 (N3899, N3885);
xor XOR2 (N3900, N3861, N364);
nand NAND2 (N3901, N3890, N299);
xor XOR2 (N3902, N3898, N2759);
or OR3 (N3903, N3899, N2342, N174);
xor XOR2 (N3904, N3903, N726);
nand NAND3 (N3905, N3894, N2218, N260);
nor NOR2 (N3906, N3897, N1888);
buf BUF1 (N3907, N3902);
nor NOR2 (N3908, N3896, N3144);
buf BUF1 (N3909, N3888);
and AND2 (N3910, N3892, N1503);
nand NAND3 (N3911, N3901, N3338, N3741);
buf BUF1 (N3912, N3907);
not NOT1 (N3913, N3905);
xor XOR2 (N3914, N3908, N410);
not NOT1 (N3915, N3900);
or OR2 (N3916, N3906, N152);
or OR4 (N3917, N3914, N3272, N62, N3466);
nand NAND2 (N3918, N3910, N1999);
or OR3 (N3919, N3917, N3208, N676);
xor XOR2 (N3920, N3916, N2597);
or OR3 (N3921, N3909, N3756, N3087);
buf BUF1 (N3922, N3904);
or OR2 (N3923, N3920, N3580);
buf BUF1 (N3924, N3922);
not NOT1 (N3925, N3912);
xor XOR2 (N3926, N3923, N1403);
or OR4 (N3927, N3924, N2472, N3909, N1796);
nor NOR4 (N3928, N3884, N1399, N7, N2927);
nand NAND4 (N3929, N3911, N1151, N807, N2213);
or OR3 (N3930, N3918, N3350, N971);
or OR3 (N3931, N3927, N2706, N1618);
buf BUF1 (N3932, N3929);
not NOT1 (N3933, N3931);
xor XOR2 (N3934, N3930, N1202);
nor NOR2 (N3935, N3928, N1004);
nor NOR2 (N3936, N3935, N2592);
and AND3 (N3937, N3921, N2919, N2468);
nor NOR3 (N3938, N3919, N2063, N3595);
buf BUF1 (N3939, N3932);
nand NAND2 (N3940, N3913, N3128);
xor XOR2 (N3941, N3926, N3529);
not NOT1 (N3942, N3933);
nand NAND2 (N3943, N3942, N2765);
or OR4 (N3944, N3937, N93, N495, N3185);
nand NAND3 (N3945, N3943, N1662, N2201);
buf BUF1 (N3946, N3938);
xor XOR2 (N3947, N3925, N3468);
buf BUF1 (N3948, N3947);
buf BUF1 (N3949, N3915);
nand NAND2 (N3950, N3941, N367);
not NOT1 (N3951, N3950);
not NOT1 (N3952, N3934);
xor XOR2 (N3953, N3944, N2448);
and AND4 (N3954, N3951, N235, N3150, N3822);
and AND2 (N3955, N3954, N2747);
nand NAND3 (N3956, N3952, N900, N3347);
and AND2 (N3957, N3939, N1100);
nor NOR3 (N3958, N3956, N1802, N1416);
not NOT1 (N3959, N3953);
buf BUF1 (N3960, N3936);
xor XOR2 (N3961, N3949, N2295);
nand NAND2 (N3962, N3960, N317);
or OR3 (N3963, N3959, N1419, N667);
nor NOR4 (N3964, N3955, N2093, N3517, N210);
buf BUF1 (N3965, N3964);
nand NAND4 (N3966, N3965, N2786, N1379, N1011);
nor NOR4 (N3967, N3940, N3439, N657, N502);
nand NAND4 (N3968, N3946, N357, N1037, N3170);
not NOT1 (N3969, N3957);
and AND3 (N3970, N3966, N761, N2920);
not NOT1 (N3971, N3945);
or OR4 (N3972, N3958, N1476, N2542, N1964);
xor XOR2 (N3973, N3969, N541);
nor NOR2 (N3974, N3967, N1127);
and AND4 (N3975, N3970, N3753, N2992, N1451);
xor XOR2 (N3976, N3972, N1931);
buf BUF1 (N3977, N3976);
nor NOR3 (N3978, N3973, N2919, N2522);
and AND4 (N3979, N3962, N1372, N448, N3928);
not NOT1 (N3980, N3978);
or OR3 (N3981, N3974, N3447, N555);
nand NAND2 (N3982, N3968, N2319);
or OR3 (N3983, N3981, N587, N319);
not NOT1 (N3984, N3963);
nor NOR2 (N3985, N3982, N209);
not NOT1 (N3986, N3948);
nand NAND4 (N3987, N3961, N2621, N1728, N143);
buf BUF1 (N3988, N3983);
not NOT1 (N3989, N3975);
and AND4 (N3990, N3985, N2656, N353, N3154);
nand NAND2 (N3991, N3977, N1540);
not NOT1 (N3992, N3984);
xor XOR2 (N3993, N3988, N2782);
buf BUF1 (N3994, N3986);
and AND2 (N3995, N3991, N3543);
and AND2 (N3996, N3989, N1374);
not NOT1 (N3997, N3994);
nor NOR4 (N3998, N3990, N3979, N2569, N663);
nand NAND4 (N3999, N165, N3093, N2038, N1921);
or OR2 (N4000, N3996, N1344);
and AND3 (N4001, N3987, N1136, N2788);
buf BUF1 (N4002, N3995);
xor XOR2 (N4003, N3997, N1570);
buf BUF1 (N4004, N4003);
nor NOR3 (N4005, N3980, N3702, N3663);
nor NOR4 (N4006, N4000, N354, N2532, N1142);
or OR2 (N4007, N4006, N2986);
or OR4 (N4008, N3992, N938, N1614, N1805);
and AND3 (N4009, N4002, N819, N2581);
or OR2 (N4010, N4009, N2456);
not NOT1 (N4011, N4007);
nand NAND2 (N4012, N3998, N1404);
not NOT1 (N4013, N3993);
nor NOR2 (N4014, N4004, N3929);
nor NOR2 (N4015, N4011, N1900);
and AND4 (N4016, N4005, N1437, N913, N2540);
buf BUF1 (N4017, N4008);
nand NAND3 (N4018, N4001, N1197, N302);
and AND3 (N4019, N4016, N2439, N339);
nor NOR2 (N4020, N4012, N3396);
and AND3 (N4021, N4010, N3670, N2423);
not NOT1 (N4022, N3999);
not NOT1 (N4023, N4018);
nor NOR2 (N4024, N3971, N523);
xor XOR2 (N4025, N4023, N3757);
nor NOR3 (N4026, N4021, N3654, N3756);
and AND2 (N4027, N4017, N2890);
and AND4 (N4028, N4026, N1703, N2900, N1820);
buf BUF1 (N4029, N4025);
nor NOR2 (N4030, N4024, N1891);
buf BUF1 (N4031, N4014);
and AND4 (N4032, N4031, N3399, N1239, N3129);
xor XOR2 (N4033, N4020, N2478);
buf BUF1 (N4034, N4030);
nor NOR4 (N4035, N4032, N130, N269, N3344);
buf BUF1 (N4036, N4029);
nand NAND2 (N4037, N4035, N3136);
and AND4 (N4038, N4015, N1647, N3547, N3573);
nor NOR3 (N4039, N4033, N1901, N3646);
buf BUF1 (N4040, N4037);
nor NOR3 (N4041, N4019, N365, N819);
nand NAND4 (N4042, N4013, N889, N2635, N2623);
xor XOR2 (N4043, N4036, N3435);
not NOT1 (N4044, N4034);
nand NAND3 (N4045, N4042, N2103, N3501);
not NOT1 (N4046, N4044);
buf BUF1 (N4047, N4039);
nand NAND4 (N4048, N4045, N1621, N347, N2515);
xor XOR2 (N4049, N4047, N47);
nand NAND3 (N4050, N4041, N295, N525);
and AND4 (N4051, N4048, N587, N3088, N1820);
xor XOR2 (N4052, N4040, N3617);
nor NOR4 (N4053, N4051, N3908, N2894, N3175);
buf BUF1 (N4054, N4053);
xor XOR2 (N4055, N4028, N3159);
and AND2 (N4056, N4038, N1332);
nor NOR3 (N4057, N4052, N3387, N3760);
nor NOR4 (N4058, N4022, N2377, N684, N1267);
nor NOR3 (N4059, N4027, N1710, N4027);
nand NAND2 (N4060, N4054, N3894);
buf BUF1 (N4061, N4060);
nor NOR3 (N4062, N4058, N3819, N1327);
or OR4 (N4063, N4059, N407, N3835, N1579);
not NOT1 (N4064, N4062);
or OR3 (N4065, N4049, N1059, N3777);
or OR3 (N4066, N4055, N2389, N2610);
or OR3 (N4067, N4056, N335, N1574);
not NOT1 (N4068, N4061);
or OR2 (N4069, N4066, N2672);
not NOT1 (N4070, N4069);
and AND3 (N4071, N4057, N2017, N1884);
or OR2 (N4072, N4071, N1926);
not NOT1 (N4073, N4065);
nor NOR3 (N4074, N4043, N3715, N3776);
nor NOR4 (N4075, N4072, N735, N1588, N2461);
nand NAND3 (N4076, N4075, N3360, N437);
xor XOR2 (N4077, N4064, N856);
and AND2 (N4078, N4074, N3983);
nor NOR3 (N4079, N4050, N3378, N1942);
nor NOR2 (N4080, N4046, N1651);
nor NOR3 (N4081, N4073, N1988, N2599);
and AND3 (N4082, N4079, N641, N2971);
xor XOR2 (N4083, N4081, N3548);
buf BUF1 (N4084, N4077);
nor NOR4 (N4085, N4076, N382, N1141, N1498);
nand NAND2 (N4086, N4063, N4051);
xor XOR2 (N4087, N4086, N500);
nand NAND2 (N4088, N4078, N3887);
not NOT1 (N4089, N4083);
xor XOR2 (N4090, N4067, N2178);
or OR2 (N4091, N4068, N3786);
nand NAND2 (N4092, N4090, N4089);
buf BUF1 (N4093, N1782);
xor XOR2 (N4094, N4084, N3085);
nor NOR3 (N4095, N4080, N3789, N682);
nor NOR4 (N4096, N4092, N1800, N3950, N2659);
nand NAND3 (N4097, N4088, N903, N632);
nor NOR4 (N4098, N4094, N3928, N1197, N860);
nor NOR4 (N4099, N4095, N1595, N1212, N296);
and AND2 (N4100, N4093, N3175);
nand NAND2 (N4101, N4100, N1609);
and AND4 (N4102, N4099, N1359, N636, N3919);
or OR3 (N4103, N4070, N2634, N928);
nand NAND4 (N4104, N4103, N1961, N1299, N2786);
or OR3 (N4105, N4098, N2273, N110);
buf BUF1 (N4106, N4102);
not NOT1 (N4107, N4104);
not NOT1 (N4108, N4082);
buf BUF1 (N4109, N4105);
xor XOR2 (N4110, N4096, N3315);
nor NOR2 (N4111, N4101, N1700);
not NOT1 (N4112, N4087);
xor XOR2 (N4113, N4106, N3974);
xor XOR2 (N4114, N4107, N115);
buf BUF1 (N4115, N4109);
and AND2 (N4116, N4113, N3180);
nand NAND3 (N4117, N4110, N3978, N338);
nand NAND3 (N4118, N4112, N2434, N1647);
nand NAND3 (N4119, N4111, N3465, N607);
xor XOR2 (N4120, N4114, N1546);
not NOT1 (N4121, N4116);
nor NOR3 (N4122, N4119, N3531, N1408);
and AND3 (N4123, N4118, N2289, N2060);
xor XOR2 (N4124, N4091, N1983);
or OR3 (N4125, N4108, N167, N894);
nor NOR3 (N4126, N4122, N1866, N2055);
nor NOR2 (N4127, N4124, N2615);
nor NOR4 (N4128, N4115, N2253, N2574, N1282);
buf BUF1 (N4129, N4121);
not NOT1 (N4130, N4085);
buf BUF1 (N4131, N4129);
nand NAND4 (N4132, N4097, N407, N1088, N3336);
nand NAND4 (N4133, N4127, N3180, N930, N804);
not NOT1 (N4134, N4125);
xor XOR2 (N4135, N4120, N2528);
xor XOR2 (N4136, N4133, N2070);
xor XOR2 (N4137, N4126, N2445);
and AND2 (N4138, N4137, N348);
buf BUF1 (N4139, N4136);
xor XOR2 (N4140, N4117, N368);
nand NAND4 (N4141, N4128, N2889, N2957, N3554);
and AND2 (N4142, N4135, N1026);
nand NAND4 (N4143, N4123, N897, N2949, N1157);
xor XOR2 (N4144, N4138, N1261);
nor NOR4 (N4145, N4134, N439, N3438, N2492);
not NOT1 (N4146, N4130);
nand NAND3 (N4147, N4141, N891, N2011);
nand NAND3 (N4148, N4144, N545, N3309);
nand NAND3 (N4149, N4131, N1750, N2567);
or OR2 (N4150, N4147, N2245);
nor NOR4 (N4151, N4143, N3222, N158, N1264);
and AND3 (N4152, N4148, N3165, N1779);
and AND2 (N4153, N4152, N2679);
xor XOR2 (N4154, N4142, N2992);
not NOT1 (N4155, N4154);
nor NOR3 (N4156, N4139, N2805, N2551);
or OR2 (N4157, N4156, N4051);
nand NAND3 (N4158, N4150, N2970, N1471);
buf BUF1 (N4159, N4157);
not NOT1 (N4160, N4158);
not NOT1 (N4161, N4151);
and AND4 (N4162, N4132, N3680, N2302, N338);
nor NOR4 (N4163, N4140, N373, N3248, N666);
buf BUF1 (N4164, N4149);
and AND2 (N4165, N4162, N3288);
and AND3 (N4166, N4155, N3155, N848);
nand NAND3 (N4167, N4165, N1797, N3702);
not NOT1 (N4168, N4161);
nand NAND4 (N4169, N4164, N3366, N1896, N3766);
buf BUF1 (N4170, N4166);
buf BUF1 (N4171, N4163);
buf BUF1 (N4172, N4159);
buf BUF1 (N4173, N4170);
xor XOR2 (N4174, N4173, N4118);
nor NOR4 (N4175, N4167, N1711, N971, N1479);
or OR3 (N4176, N4153, N1543, N3905);
not NOT1 (N4177, N4171);
or OR4 (N4178, N4168, N1418, N3347, N2513);
not NOT1 (N4179, N4172);
not NOT1 (N4180, N4177);
and AND4 (N4181, N4180, N180, N37, N2430);
xor XOR2 (N4182, N4176, N3167);
or OR4 (N4183, N4145, N3602, N294, N3641);
xor XOR2 (N4184, N4174, N467);
nor NOR3 (N4185, N4146, N3707, N882);
xor XOR2 (N4186, N4183, N735);
xor XOR2 (N4187, N4175, N3236);
nor NOR4 (N4188, N4182, N2310, N2112, N1318);
and AND2 (N4189, N4185, N1510);
buf BUF1 (N4190, N4181);
nand NAND2 (N4191, N4178, N3543);
buf BUF1 (N4192, N4189);
not NOT1 (N4193, N4192);
and AND3 (N4194, N4190, N1127, N630);
and AND2 (N4195, N4169, N1165);
and AND4 (N4196, N4187, N1032, N444, N2922);
buf BUF1 (N4197, N4194);
nor NOR3 (N4198, N4179, N2687, N1666);
xor XOR2 (N4199, N4195, N1467);
nand NAND3 (N4200, N4186, N596, N1981);
and AND4 (N4201, N4197, N804, N3605, N3663);
not NOT1 (N4202, N4201);
not NOT1 (N4203, N4160);
nor NOR3 (N4204, N4200, N3657, N3268);
nand NAND2 (N4205, N4188, N3020);
nand NAND4 (N4206, N4203, N600, N550, N1330);
or OR4 (N4207, N4198, N983, N319, N4037);
buf BUF1 (N4208, N4199);
and AND4 (N4209, N4208, N3936, N2568, N2550);
or OR4 (N4210, N4193, N988, N3422, N1428);
or OR4 (N4211, N4206, N2005, N1414, N2933);
xor XOR2 (N4212, N4196, N3971);
not NOT1 (N4213, N4205);
buf BUF1 (N4214, N4210);
not NOT1 (N4215, N4213);
not NOT1 (N4216, N4207);
nand NAND2 (N4217, N4211, N907);
nor NOR3 (N4218, N4204, N1038, N4003);
nor NOR4 (N4219, N4191, N3423, N3886, N1777);
or OR4 (N4220, N4184, N641, N3480, N3474);
or OR4 (N4221, N4215, N2426, N3256, N3943);
buf BUF1 (N4222, N4214);
not NOT1 (N4223, N4222);
not NOT1 (N4224, N4220);
nor NOR4 (N4225, N4216, N79, N3840, N2976);
and AND3 (N4226, N4218, N413, N3433);
xor XOR2 (N4227, N4202, N359);
buf BUF1 (N4228, N4225);
nor NOR3 (N4229, N4219, N2285, N3661);
and AND3 (N4230, N4209, N1538, N2778);
xor XOR2 (N4231, N4221, N4172);
nor NOR3 (N4232, N4223, N718, N233);
nand NAND3 (N4233, N4228, N758, N2313);
xor XOR2 (N4234, N4224, N4059);
buf BUF1 (N4235, N4226);
or OR4 (N4236, N4232, N49, N4049, N1356);
buf BUF1 (N4237, N4217);
or OR4 (N4238, N4230, N4235, N421, N3358);
buf BUF1 (N4239, N2966);
nor NOR3 (N4240, N4239, N663, N1245);
xor XOR2 (N4241, N4240, N2645);
nor NOR4 (N4242, N4236, N2129, N3440, N1728);
nor NOR2 (N4243, N4233, N382);
or OR2 (N4244, N4234, N3056);
nand NAND4 (N4245, N4243, N4174, N2747, N3869);
nor NOR3 (N4246, N4245, N2465, N2739);
nand NAND3 (N4247, N4244, N2955, N2483);
xor XOR2 (N4248, N4227, N312);
and AND2 (N4249, N4212, N3877);
nor NOR3 (N4250, N4249, N3080, N4038);
nand NAND4 (N4251, N4241, N2360, N3032, N55);
not NOT1 (N4252, N4237);
xor XOR2 (N4253, N4252, N430);
or OR3 (N4254, N4251, N637, N907);
and AND4 (N4255, N4229, N1399, N2185, N3404);
not NOT1 (N4256, N4255);
or OR3 (N4257, N4248, N1566, N698);
buf BUF1 (N4258, N4231);
and AND2 (N4259, N4247, N730);
xor XOR2 (N4260, N4250, N2036);
buf BUF1 (N4261, N4238);
xor XOR2 (N4262, N4256, N772);
nor NOR2 (N4263, N4259, N1146);
or OR3 (N4264, N4262, N3897, N3086);
and AND2 (N4265, N4260, N3784);
nand NAND4 (N4266, N4261, N1590, N2096, N198);
and AND2 (N4267, N4263, N683);
xor XOR2 (N4268, N4242, N3203);
nand NAND4 (N4269, N4246, N2403, N943, N2592);
buf BUF1 (N4270, N4253);
and AND3 (N4271, N4269, N4153, N1502);
not NOT1 (N4272, N4257);
nor NOR4 (N4273, N4272, N1934, N1304, N2570);
and AND2 (N4274, N4264, N2422);
and AND4 (N4275, N4270, N3864, N1025, N1622);
xor XOR2 (N4276, N4274, N2793);
and AND3 (N4277, N4273, N2877, N3354);
buf BUF1 (N4278, N4266);
xor XOR2 (N4279, N4278, N4199);
and AND2 (N4280, N4279, N919);
not NOT1 (N4281, N4267);
not NOT1 (N4282, N4276);
and AND4 (N4283, N4282, N4169, N619, N2268);
and AND2 (N4284, N4254, N789);
xor XOR2 (N4285, N4284, N267);
and AND3 (N4286, N4285, N1849, N4132);
or OR4 (N4287, N4271, N803, N1034, N452);
or OR2 (N4288, N4277, N4202);
nand NAND2 (N4289, N4281, N1936);
not NOT1 (N4290, N4268);
nand NAND2 (N4291, N4280, N3417);
or OR2 (N4292, N4286, N175);
or OR3 (N4293, N4275, N1632, N1443);
buf BUF1 (N4294, N4265);
buf BUF1 (N4295, N4294);
not NOT1 (N4296, N4258);
and AND2 (N4297, N4283, N1098);
xor XOR2 (N4298, N4288, N1726);
nand NAND4 (N4299, N4291, N729, N972, N75);
buf BUF1 (N4300, N4293);
or OR4 (N4301, N4296, N4115, N325, N2211);
buf BUF1 (N4302, N4297);
nand NAND3 (N4303, N4301, N1994, N36);
xor XOR2 (N4304, N4302, N3216);
not NOT1 (N4305, N4290);
nand NAND3 (N4306, N4289, N4203, N2530);
buf BUF1 (N4307, N4287);
not NOT1 (N4308, N4295);
or OR3 (N4309, N4304, N2843, N3252);
nor NOR3 (N4310, N4309, N1567, N1312);
xor XOR2 (N4311, N4300, N2699);
nor NOR4 (N4312, N4307, N726, N3989, N1371);
xor XOR2 (N4313, N4303, N3137);
nor NOR3 (N4314, N4299, N3107, N3139);
and AND4 (N4315, N4298, N1906, N167, N2971);
and AND2 (N4316, N4315, N3723);
nand NAND4 (N4317, N4316, N489, N3500, N3645);
nand NAND3 (N4318, N4311, N1321, N2669);
not NOT1 (N4319, N4292);
xor XOR2 (N4320, N4312, N2566);
nand NAND3 (N4321, N4318, N1180, N3828);
buf BUF1 (N4322, N4320);
nor NOR2 (N4323, N4322, N3564);
not NOT1 (N4324, N4319);
nand NAND4 (N4325, N4314, N1464, N3279, N3960);
xor XOR2 (N4326, N4321, N2158);
not NOT1 (N4327, N4306);
nor NOR4 (N4328, N4323, N818, N868, N2228);
xor XOR2 (N4329, N4326, N1703);
xor XOR2 (N4330, N4328, N1398);
nor NOR3 (N4331, N4313, N1690, N2948);
nor NOR2 (N4332, N4305, N2737);
nand NAND2 (N4333, N4324, N2634);
buf BUF1 (N4334, N4330);
buf BUF1 (N4335, N4334);
nor NOR3 (N4336, N4325, N3767, N1489);
xor XOR2 (N4337, N4329, N1306);
or OR3 (N4338, N4331, N3755, N2021);
not NOT1 (N4339, N4337);
xor XOR2 (N4340, N4327, N2548);
nor NOR4 (N4341, N4317, N1452, N811, N459);
nand NAND2 (N4342, N4338, N3056);
and AND4 (N4343, N4342, N4062, N353, N2755);
buf BUF1 (N4344, N4339);
not NOT1 (N4345, N4308);
nand NAND2 (N4346, N4344, N253);
nand NAND3 (N4347, N4335, N2178, N2528);
not NOT1 (N4348, N4346);
nand NAND2 (N4349, N4347, N3251);
and AND4 (N4350, N4332, N2889, N205, N2385);
nor NOR3 (N4351, N4310, N1037, N1079);
not NOT1 (N4352, N4336);
nand NAND3 (N4353, N4349, N2724, N1129);
nor NOR4 (N4354, N4353, N1090, N2629, N3487);
not NOT1 (N4355, N4351);
or OR2 (N4356, N4341, N311);
and AND4 (N4357, N4345, N2995, N2045, N3760);
nor NOR4 (N4358, N4348, N323, N1387, N1014);
not NOT1 (N4359, N4357);
buf BUF1 (N4360, N4352);
or OR4 (N4361, N4343, N1228, N1446, N482);
xor XOR2 (N4362, N4354, N944);
xor XOR2 (N4363, N4350, N1307);
and AND4 (N4364, N4361, N1829, N2178, N3283);
nand NAND4 (N4365, N4356, N2069, N2601, N3941);
nor NOR2 (N4366, N4355, N2861);
or OR2 (N4367, N4366, N1251);
xor XOR2 (N4368, N4362, N303);
nand NAND4 (N4369, N4360, N912, N2691, N966);
and AND4 (N4370, N4363, N4085, N1841, N3463);
and AND2 (N4371, N4364, N1242);
and AND4 (N4372, N4371, N4329, N2877, N2710);
nor NOR2 (N4373, N4370, N1217);
buf BUF1 (N4374, N4368);
not NOT1 (N4375, N4359);
not NOT1 (N4376, N4333);
xor XOR2 (N4377, N4367, N2661);
xor XOR2 (N4378, N4375, N338);
buf BUF1 (N4379, N4373);
nor NOR4 (N4380, N4379, N3747, N4336, N1975);
nand NAND3 (N4381, N4365, N152, N109);
not NOT1 (N4382, N4381);
xor XOR2 (N4383, N4378, N2054);
and AND2 (N4384, N4374, N202);
xor XOR2 (N4385, N4383, N3509);
nor NOR4 (N4386, N4340, N2252, N24, N3099);
nor NOR3 (N4387, N4384, N2607, N3938);
buf BUF1 (N4388, N4369);
buf BUF1 (N4389, N4358);
and AND4 (N4390, N4385, N4338, N2672, N1270);
nand NAND3 (N4391, N4376, N3182, N3367);
and AND3 (N4392, N4382, N4073, N2398);
and AND4 (N4393, N4386, N992, N343, N3966);
nor NOR3 (N4394, N4387, N2740, N3826);
buf BUF1 (N4395, N4377);
nor NOR2 (N4396, N4395, N1144);
not NOT1 (N4397, N4391);
xor XOR2 (N4398, N4390, N975);
not NOT1 (N4399, N4393);
not NOT1 (N4400, N4388);
nand NAND2 (N4401, N4398, N1172);
not NOT1 (N4402, N4399);
nor NOR3 (N4403, N4402, N512, N135);
xor XOR2 (N4404, N4396, N1645);
not NOT1 (N4405, N4394);
or OR3 (N4406, N4397, N4269, N3097);
not NOT1 (N4407, N4403);
or OR2 (N4408, N4407, N934);
buf BUF1 (N4409, N4408);
nor NOR4 (N4410, N4405, N2508, N1353, N1046);
buf BUF1 (N4411, N4404);
nand NAND2 (N4412, N4401, N3381);
buf BUF1 (N4413, N4412);
buf BUF1 (N4414, N4410);
and AND2 (N4415, N4409, N3439);
not NOT1 (N4416, N4415);
nand NAND4 (N4417, N4392, N1433, N3054, N1330);
or OR2 (N4418, N4414, N3746);
buf BUF1 (N4419, N4413);
and AND3 (N4420, N4400, N2732, N2834);
buf BUF1 (N4421, N4372);
buf BUF1 (N4422, N4416);
and AND3 (N4423, N4418, N2909, N120);
nand NAND4 (N4424, N4420, N1931, N2361, N3817);
buf BUF1 (N4425, N4417);
buf BUF1 (N4426, N4389);
xor XOR2 (N4427, N4425, N3272);
nor NOR4 (N4428, N4380, N2143, N1985, N3843);
nor NOR3 (N4429, N4422, N2987, N2301);
nor NOR2 (N4430, N4429, N2166);
or OR4 (N4431, N4411, N2786, N495, N1574);
and AND2 (N4432, N4421, N2859);
nor NOR2 (N4433, N4427, N4047);
nor NOR3 (N4434, N4428, N3444, N643);
not NOT1 (N4435, N4433);
or OR2 (N4436, N4423, N361);
and AND4 (N4437, N4430, N1349, N1626, N2241);
and AND2 (N4438, N4424, N1545);
and AND3 (N4439, N4431, N1540, N2932);
nor NOR2 (N4440, N4406, N1816);
or OR2 (N4441, N4434, N1577);
or OR3 (N4442, N4419, N3630, N2710);
not NOT1 (N4443, N4436);
not NOT1 (N4444, N4441);
not NOT1 (N4445, N4443);
nor NOR2 (N4446, N4444, N987);
not NOT1 (N4447, N4442);
not NOT1 (N4448, N4438);
nand NAND2 (N4449, N4440, N215);
buf BUF1 (N4450, N4445);
buf BUF1 (N4451, N4432);
and AND4 (N4452, N4435, N755, N941, N4132);
xor XOR2 (N4453, N4426, N2002);
xor XOR2 (N4454, N4451, N3018);
xor XOR2 (N4455, N4439, N2525);
nor NOR3 (N4456, N4437, N3147, N4267);
and AND2 (N4457, N4447, N4349);
not NOT1 (N4458, N4454);
nand NAND2 (N4459, N4457, N4447);
nor NOR4 (N4460, N4455, N255, N4412, N2947);
buf BUF1 (N4461, N4459);
not NOT1 (N4462, N4458);
nand NAND2 (N4463, N4450, N2249);
nand NAND4 (N4464, N4461, N1386, N442, N269);
nand NAND2 (N4465, N4448, N2853);
xor XOR2 (N4466, N4452, N2654);
nor NOR4 (N4467, N4460, N2145, N1039, N1181);
and AND2 (N4468, N4462, N3152);
not NOT1 (N4469, N4464);
nand NAND3 (N4470, N4469, N3411, N2147);
nor NOR4 (N4471, N4468, N2869, N1706, N747);
nand NAND4 (N4472, N4470, N2653, N2472, N143);
nand NAND4 (N4473, N4471, N1795, N3583, N1555);
or OR4 (N4474, N4449, N1135, N3128, N1373);
nor NOR3 (N4475, N4446, N3082, N688);
xor XOR2 (N4476, N4463, N1488);
not NOT1 (N4477, N4473);
nor NOR3 (N4478, N4476, N1765, N1058);
xor XOR2 (N4479, N4478, N3794);
not NOT1 (N4480, N4475);
or OR4 (N4481, N4477, N3705, N3956, N2030);
not NOT1 (N4482, N4465);
and AND4 (N4483, N4472, N2924, N2433, N948);
nor NOR3 (N4484, N4483, N4399, N594);
buf BUF1 (N4485, N4467);
nand NAND2 (N4486, N4481, N1318);
and AND2 (N4487, N4486, N2362);
nand NAND3 (N4488, N4485, N1909, N4252);
or OR3 (N4489, N4484, N500, N3408);
nor NOR4 (N4490, N4482, N2416, N732, N3045);
or OR2 (N4491, N4487, N3968);
buf BUF1 (N4492, N4466);
nand NAND2 (N4493, N4453, N3557);
nor NOR4 (N4494, N4488, N334, N2077, N1377);
nand NAND2 (N4495, N4493, N3236);
nor NOR3 (N4496, N4491, N2573, N897);
not NOT1 (N4497, N4490);
or OR3 (N4498, N4480, N4394, N2983);
not NOT1 (N4499, N4498);
not NOT1 (N4500, N4499);
and AND2 (N4501, N4492, N4107);
not NOT1 (N4502, N4489);
or OR3 (N4503, N4497, N1208, N3743);
nor NOR2 (N4504, N4479, N290);
buf BUF1 (N4505, N4494);
or OR2 (N4506, N4504, N2096);
xor XOR2 (N4507, N4502, N2547);
or OR3 (N4508, N4507, N2748, N2997);
buf BUF1 (N4509, N4495);
and AND4 (N4510, N4508, N1774, N745, N623);
xor XOR2 (N4511, N4496, N4377);
buf BUF1 (N4512, N4510);
buf BUF1 (N4513, N4503);
nor NOR4 (N4514, N4513, N135, N889, N912);
or OR3 (N4515, N4474, N2734, N537);
not NOT1 (N4516, N4511);
and AND3 (N4517, N4500, N4476, N969);
or OR2 (N4518, N4514, N605);
nand NAND2 (N4519, N4512, N3876);
and AND3 (N4520, N4515, N3450, N3462);
nor NOR3 (N4521, N4517, N2371, N3169);
xor XOR2 (N4522, N4456, N791);
nand NAND4 (N4523, N4509, N4252, N3531, N3119);
or OR4 (N4524, N4523, N3389, N2590, N648);
not NOT1 (N4525, N4501);
not NOT1 (N4526, N4524);
and AND2 (N4527, N4516, N2115);
nand NAND4 (N4528, N4527, N4114, N3601, N517);
xor XOR2 (N4529, N4505, N2156);
xor XOR2 (N4530, N4526, N605);
buf BUF1 (N4531, N4518);
nand NAND3 (N4532, N4528, N1086, N3684);
and AND2 (N4533, N4519, N607);
xor XOR2 (N4534, N4521, N2358);
buf BUF1 (N4535, N4532);
and AND3 (N4536, N4534, N1194, N3601);
nor NOR4 (N4537, N4522, N3618, N3542, N66);
not NOT1 (N4538, N4520);
buf BUF1 (N4539, N4530);
nor NOR2 (N4540, N4537, N1389);
and AND3 (N4541, N4531, N3751, N3160);
nor NOR4 (N4542, N4535, N882, N2658, N465);
xor XOR2 (N4543, N4525, N4254);
xor XOR2 (N4544, N4533, N2175);
and AND4 (N4545, N4543, N425, N2612, N2686);
nand NAND3 (N4546, N4538, N3696, N107);
nor NOR4 (N4547, N4546, N4359, N1979, N3061);
nor NOR4 (N4548, N4506, N3303, N1393, N2498);
nand NAND2 (N4549, N4536, N1582);
not NOT1 (N4550, N4544);
nor NOR3 (N4551, N4549, N3389, N286);
nand NAND4 (N4552, N4541, N45, N2450, N518);
or OR3 (N4553, N4529, N3230, N2483);
xor XOR2 (N4554, N4540, N3966);
nand NAND3 (N4555, N4551, N551, N2036);
buf BUF1 (N4556, N4548);
xor XOR2 (N4557, N4550, N113);
not NOT1 (N4558, N4553);
or OR4 (N4559, N4547, N1579, N4089, N399);
not NOT1 (N4560, N4545);
xor XOR2 (N4561, N4558, N4221);
nand NAND3 (N4562, N4539, N2812, N3243);
not NOT1 (N4563, N4552);
nor NOR4 (N4564, N4556, N1745, N2822, N396);
or OR2 (N4565, N4554, N2800);
buf BUF1 (N4566, N4561);
and AND2 (N4567, N4565, N2308);
nand NAND2 (N4568, N4542, N3253);
not NOT1 (N4569, N4566);
nand NAND4 (N4570, N4562, N2595, N542, N1132);
or OR3 (N4571, N4557, N3528, N3962);
and AND4 (N4572, N4569, N1172, N2178, N389);
nor NOR2 (N4573, N4572, N608);
and AND2 (N4574, N4559, N4520);
buf BUF1 (N4575, N4571);
and AND4 (N4576, N4570, N1386, N116, N500);
xor XOR2 (N4577, N4560, N4492);
not NOT1 (N4578, N4576);
xor XOR2 (N4579, N4573, N1437);
nor NOR2 (N4580, N4563, N3832);
or OR4 (N4581, N4568, N4456, N1300, N2731);
or OR2 (N4582, N4574, N2724);
not NOT1 (N4583, N4575);
and AND3 (N4584, N4579, N2964, N1135);
or OR3 (N4585, N4578, N376, N785);
nor NOR2 (N4586, N4555, N1623);
not NOT1 (N4587, N4564);
xor XOR2 (N4588, N4577, N1348);
nor NOR2 (N4589, N4585, N2449);
nor NOR4 (N4590, N4567, N1145, N132, N2402);
nand NAND3 (N4591, N4588, N1659, N3197);
nor NOR2 (N4592, N4581, N518);
nand NAND2 (N4593, N4582, N4061);
nor NOR3 (N4594, N4590, N965, N1005);
nor NOR2 (N4595, N4592, N4185);
not NOT1 (N4596, N4595);
xor XOR2 (N4597, N4586, N1730);
not NOT1 (N4598, N4587);
xor XOR2 (N4599, N4584, N3196);
nand NAND3 (N4600, N4583, N4206, N2772);
xor XOR2 (N4601, N4600, N898);
not NOT1 (N4602, N4580);
xor XOR2 (N4603, N4602, N4373);
not NOT1 (N4604, N4589);
nand NAND3 (N4605, N4598, N4312, N1445);
xor XOR2 (N4606, N4603, N1104);
and AND3 (N4607, N4593, N4123, N3552);
or OR3 (N4608, N4601, N2338, N45);
or OR2 (N4609, N4594, N3695);
nand NAND4 (N4610, N4591, N2754, N156, N2607);
or OR3 (N4611, N4606, N2271, N4346);
nor NOR3 (N4612, N4611, N3470, N4325);
nand NAND4 (N4613, N4599, N2263, N2647, N3165);
not NOT1 (N4614, N4608);
not NOT1 (N4615, N4614);
or OR3 (N4616, N4607, N4291, N2559);
not NOT1 (N4617, N4615);
xor XOR2 (N4618, N4596, N4160);
or OR2 (N4619, N4617, N2357);
or OR2 (N4620, N4618, N4200);
or OR3 (N4621, N4616, N1734, N3492);
xor XOR2 (N4622, N4604, N3861);
xor XOR2 (N4623, N4597, N3168);
buf BUF1 (N4624, N4612);
not NOT1 (N4625, N4620);
nor NOR2 (N4626, N4623, N2508);
not NOT1 (N4627, N4613);
nand NAND3 (N4628, N4627, N4416, N30);
not NOT1 (N4629, N4622);
or OR4 (N4630, N4628, N980, N168, N1212);
nor NOR4 (N4631, N4625, N518, N377, N2484);
not NOT1 (N4632, N4610);
buf BUF1 (N4633, N4624);
nor NOR4 (N4634, N4631, N1127, N3801, N4316);
buf BUF1 (N4635, N4605);
nor NOR3 (N4636, N4626, N1777, N222);
buf BUF1 (N4637, N4635);
nand NAND3 (N4638, N4633, N316, N3584);
nand NAND4 (N4639, N4619, N1182, N1243, N3804);
buf BUF1 (N4640, N4636);
not NOT1 (N4641, N4637);
not NOT1 (N4642, N4638);
nand NAND2 (N4643, N4621, N574);
not NOT1 (N4644, N4632);
not NOT1 (N4645, N4634);
xor XOR2 (N4646, N4609, N1328);
not NOT1 (N4647, N4641);
and AND4 (N4648, N4646, N173, N536, N1504);
or OR3 (N4649, N4630, N230, N1210);
xor XOR2 (N4650, N4642, N3273);
or OR4 (N4651, N4643, N4593, N914, N732);
nand NAND4 (N4652, N4629, N1695, N4077, N4062);
xor XOR2 (N4653, N4639, N2103);
xor XOR2 (N4654, N4647, N240);
or OR2 (N4655, N4645, N2141);
nor NOR2 (N4656, N4648, N2406);
not NOT1 (N4657, N4653);
nor NOR3 (N4658, N4654, N4458, N4226);
buf BUF1 (N4659, N4651);
not NOT1 (N4660, N4649);
xor XOR2 (N4661, N4644, N2707);
and AND4 (N4662, N4656, N3573, N147, N3221);
xor XOR2 (N4663, N4640, N4604);
xor XOR2 (N4664, N4652, N1045);
not NOT1 (N4665, N4657);
nand NAND3 (N4666, N4659, N2062, N2007);
nand NAND3 (N4667, N4650, N2280, N1346);
nor NOR2 (N4668, N4661, N2914);
xor XOR2 (N4669, N4666, N2994);
or OR3 (N4670, N4667, N2203, N820);
or OR2 (N4671, N4669, N916);
buf BUF1 (N4672, N4658);
nor NOR3 (N4673, N4671, N2083, N2438);
nand NAND3 (N4674, N4662, N3504, N83);
not NOT1 (N4675, N4663);
nand NAND2 (N4676, N4672, N1683);
or OR4 (N4677, N4665, N1788, N1908, N3587);
xor XOR2 (N4678, N4677, N79);
nor NOR4 (N4679, N4675, N4124, N3512, N15);
or OR2 (N4680, N4660, N3105);
xor XOR2 (N4681, N4674, N2035);
buf BUF1 (N4682, N4680);
and AND4 (N4683, N4664, N4650, N4529, N1217);
nor NOR3 (N4684, N4676, N1649, N1078);
not NOT1 (N4685, N4684);
nand NAND2 (N4686, N4685, N538);
buf BUF1 (N4687, N4686);
and AND2 (N4688, N4682, N3879);
buf BUF1 (N4689, N4670);
buf BUF1 (N4690, N4683);
xor XOR2 (N4691, N4668, N282);
not NOT1 (N4692, N4678);
and AND4 (N4693, N4687, N4442, N687, N3674);
not NOT1 (N4694, N4688);
nor NOR2 (N4695, N4690, N1980);
not NOT1 (N4696, N4679);
buf BUF1 (N4697, N4694);
and AND2 (N4698, N4695, N966);
or OR4 (N4699, N4696, N3948, N3651, N3579);
xor XOR2 (N4700, N4692, N145);
xor XOR2 (N4701, N4700, N1291);
and AND4 (N4702, N4697, N1855, N1667, N3216);
and AND3 (N4703, N4691, N2654, N3197);
or OR3 (N4704, N4673, N2410, N2591);
nand NAND2 (N4705, N4703, N211);
xor XOR2 (N4706, N4693, N1078);
not NOT1 (N4707, N4689);
xor XOR2 (N4708, N4699, N1989);
xor XOR2 (N4709, N4705, N1067);
not NOT1 (N4710, N4681);
nor NOR3 (N4711, N4706, N754, N1829);
nor NOR4 (N4712, N4711, N2451, N2520, N4464);
buf BUF1 (N4713, N4698);
nand NAND3 (N4714, N4708, N756, N770);
buf BUF1 (N4715, N4701);
and AND2 (N4716, N4702, N1771);
or OR3 (N4717, N4704, N1164, N3854);
nor NOR2 (N4718, N4655, N3405);
not NOT1 (N4719, N4707);
not NOT1 (N4720, N4713);
nand NAND3 (N4721, N4717, N1748, N118);
not NOT1 (N4722, N4716);
or OR2 (N4723, N4722, N2841);
buf BUF1 (N4724, N4723);
and AND4 (N4725, N4718, N3950, N4220, N147);
xor XOR2 (N4726, N4724, N2885);
or OR4 (N4727, N4726, N3932, N3349, N3116);
not NOT1 (N4728, N4712);
nand NAND3 (N4729, N4709, N2973, N3360);
or OR3 (N4730, N4729, N945, N4165);
nor NOR4 (N4731, N4721, N4080, N2478, N3074);
and AND3 (N4732, N4725, N962, N2356);
nor NOR3 (N4733, N4731, N667, N4705);
xor XOR2 (N4734, N4714, N2821);
xor XOR2 (N4735, N4727, N969);
xor XOR2 (N4736, N4732, N882);
nand NAND4 (N4737, N4735, N1403, N4526, N454);
not NOT1 (N4738, N4736);
or OR4 (N4739, N4738, N1437, N4206, N1626);
or OR3 (N4740, N4728, N4220, N3769);
or OR3 (N4741, N4734, N120, N2685);
nand NAND3 (N4742, N4741, N307, N4045);
nand NAND2 (N4743, N4740, N293);
not NOT1 (N4744, N4733);
and AND4 (N4745, N4730, N4147, N1981, N4180);
or OR4 (N4746, N4743, N3458, N1604, N4561);
xor XOR2 (N4747, N4742, N3560);
nand NAND2 (N4748, N4710, N1662);
nand NAND3 (N4749, N4748, N3642, N782);
buf BUF1 (N4750, N4749);
or OR3 (N4751, N4750, N2929, N1170);
buf BUF1 (N4752, N4719);
and AND2 (N4753, N4745, N2907);
nand NAND4 (N4754, N4737, N304, N635, N2421);
buf BUF1 (N4755, N4754);
and AND2 (N4756, N4752, N1192);
xor XOR2 (N4757, N4720, N2098);
or OR3 (N4758, N4753, N3597, N2841);
or OR4 (N4759, N4746, N4119, N191, N4643);
xor XOR2 (N4760, N4739, N1294);
or OR3 (N4761, N4760, N1012, N1936);
or OR2 (N4762, N4758, N1583);
buf BUF1 (N4763, N4755);
buf BUF1 (N4764, N4762);
nor NOR2 (N4765, N4757, N4011);
xor XOR2 (N4766, N4751, N3714);
nor NOR3 (N4767, N4763, N979, N1840);
nor NOR4 (N4768, N4759, N2553, N2482, N3490);
xor XOR2 (N4769, N4767, N2048);
nor NOR3 (N4770, N4766, N1864, N1121);
buf BUF1 (N4771, N4769);
nor NOR3 (N4772, N4715, N868, N4055);
nand NAND3 (N4773, N4768, N3721, N1342);
nor NOR4 (N4774, N4744, N2717, N297, N3707);
and AND2 (N4775, N4771, N104);
buf BUF1 (N4776, N4773);
xor XOR2 (N4777, N4770, N3874);
or OR2 (N4778, N4765, N1935);
nand NAND2 (N4779, N4747, N2059);
and AND2 (N4780, N4772, N4673);
nand NAND3 (N4781, N4779, N1911, N2893);
xor XOR2 (N4782, N4780, N3361);
nand NAND2 (N4783, N4756, N967);
nor NOR4 (N4784, N4764, N897, N3769, N2308);
xor XOR2 (N4785, N4777, N1583);
nand NAND4 (N4786, N4778, N3345, N161, N4752);
nand NAND4 (N4787, N4774, N3456, N3966, N2394);
or OR2 (N4788, N4785, N4283);
or OR3 (N4789, N4776, N2622, N1623);
nor NOR3 (N4790, N4761, N1033, N269);
or OR3 (N4791, N4788, N3988, N1947);
xor XOR2 (N4792, N4775, N865);
nor NOR2 (N4793, N4783, N3980);
not NOT1 (N4794, N4784);
nand NAND2 (N4795, N4786, N3376);
xor XOR2 (N4796, N4795, N1035);
not NOT1 (N4797, N4781);
nor NOR4 (N4798, N4797, N3321, N664, N4262);
xor XOR2 (N4799, N4782, N2830);
nand NAND2 (N4800, N4793, N2071);
nor NOR3 (N4801, N4798, N2144, N1075);
nor NOR2 (N4802, N4796, N3098);
not NOT1 (N4803, N4792);
nand NAND4 (N4804, N4787, N4550, N1860, N1286);
not NOT1 (N4805, N4803);
xor XOR2 (N4806, N4801, N3413);
buf BUF1 (N4807, N4790);
buf BUF1 (N4808, N4800);
and AND4 (N4809, N4794, N1029, N4604, N2470);
and AND2 (N4810, N4808, N726);
xor XOR2 (N4811, N4805, N360);
xor XOR2 (N4812, N4799, N3527);
not NOT1 (N4813, N4811);
nor NOR2 (N4814, N4807, N3819);
and AND3 (N4815, N4810, N1278, N2469);
nand NAND3 (N4816, N4815, N1487, N410);
xor XOR2 (N4817, N4814, N3584);
and AND2 (N4818, N4789, N4061);
nand NAND2 (N4819, N4813, N4719);
or OR4 (N4820, N4806, N4800, N4781, N2567);
not NOT1 (N4821, N4809);
or OR2 (N4822, N4820, N1043);
buf BUF1 (N4823, N4819);
buf BUF1 (N4824, N4804);
and AND4 (N4825, N4802, N2800, N3361, N2213);
nor NOR3 (N4826, N4818, N1636, N3929);
nand NAND2 (N4827, N4791, N200);
or OR4 (N4828, N4816, N3738, N3631, N2882);
or OR2 (N4829, N4824, N1229);
nand NAND2 (N4830, N4829, N1696);
nand NAND4 (N4831, N4817, N611, N1510, N2368);
xor XOR2 (N4832, N4831, N3572);
and AND4 (N4833, N4830, N4743, N1518, N640);
not NOT1 (N4834, N4821);
nor NOR3 (N4835, N4823, N359, N3358);
xor XOR2 (N4836, N4833, N2701);
buf BUF1 (N4837, N4834);
nand NAND4 (N4838, N4836, N3175, N2215, N3753);
nor NOR2 (N4839, N4832, N4675);
xor XOR2 (N4840, N4828, N4212);
or OR2 (N4841, N4839, N708);
buf BUF1 (N4842, N4840);
buf BUF1 (N4843, N4822);
not NOT1 (N4844, N4838);
not NOT1 (N4845, N4826);
or OR2 (N4846, N4844, N1359);
not NOT1 (N4847, N4842);
xor XOR2 (N4848, N4827, N1948);
xor XOR2 (N4849, N4841, N3542);
nor NOR4 (N4850, N4837, N1389, N2988, N3900);
xor XOR2 (N4851, N4848, N476);
or OR3 (N4852, N4825, N3881, N4015);
xor XOR2 (N4853, N4851, N668);
xor XOR2 (N4854, N4847, N3372);
or OR2 (N4855, N4812, N4732);
nor NOR3 (N4856, N4852, N1156, N2972);
and AND4 (N4857, N4835, N3400, N2322, N1824);
nand NAND3 (N4858, N4854, N3586, N487);
xor XOR2 (N4859, N4856, N4809);
xor XOR2 (N4860, N4859, N2988);
buf BUF1 (N4861, N4858);
xor XOR2 (N4862, N4861, N1131);
xor XOR2 (N4863, N4849, N3434);
not NOT1 (N4864, N4860);
buf BUF1 (N4865, N4843);
not NOT1 (N4866, N4864);
or OR2 (N4867, N4857, N2992);
nor NOR2 (N4868, N4862, N2660);
nor NOR2 (N4869, N4866, N2441);
buf BUF1 (N4870, N4853);
xor XOR2 (N4871, N4855, N4619);
xor XOR2 (N4872, N4863, N4713);
or OR2 (N4873, N4871, N2572);
nor NOR3 (N4874, N4846, N2735, N4382);
and AND4 (N4875, N4869, N2142, N2154, N1389);
and AND2 (N4876, N4850, N871);
or OR4 (N4877, N4870, N2267, N2564, N1105);
buf BUF1 (N4878, N4872);
or OR2 (N4879, N4876, N4106);
xor XOR2 (N4880, N4868, N2808);
nor NOR2 (N4881, N4879, N1243);
or OR4 (N4882, N4865, N2960, N1620, N2644);
and AND4 (N4883, N4881, N2588, N724, N3600);
and AND4 (N4884, N4873, N3948, N1632, N4174);
xor XOR2 (N4885, N4882, N1945);
or OR2 (N4886, N4883, N4300);
nand NAND2 (N4887, N4884, N3163);
or OR3 (N4888, N4874, N3968, N2956);
xor XOR2 (N4889, N4888, N1136);
xor XOR2 (N4890, N4880, N3300);
not NOT1 (N4891, N4886);
nand NAND4 (N4892, N4878, N1895, N1290, N1461);
xor XOR2 (N4893, N4889, N3258);
nand NAND3 (N4894, N4877, N1663, N2174);
not NOT1 (N4895, N4867);
nor NOR4 (N4896, N4892, N3682, N3607, N3716);
nand NAND3 (N4897, N4890, N3104, N4081);
or OR3 (N4898, N4893, N408, N1536);
or OR2 (N4899, N4896, N2958);
nand NAND4 (N4900, N4875, N2058, N1919, N3276);
nand NAND3 (N4901, N4845, N4502, N2235);
not NOT1 (N4902, N4900);
xor XOR2 (N4903, N4891, N725);
and AND4 (N4904, N4899, N3719, N2821, N1691);
xor XOR2 (N4905, N4887, N3021);
nor NOR2 (N4906, N4897, N244);
buf BUF1 (N4907, N4906);
nand NAND4 (N4908, N4902, N2934, N1860, N3301);
or OR4 (N4909, N4898, N1453, N2600, N4653);
or OR4 (N4910, N4904, N538, N3298, N4862);
and AND3 (N4911, N4885, N2630, N2318);
or OR3 (N4912, N4909, N1314, N2294);
nor NOR2 (N4913, N4895, N3088);
nand NAND2 (N4914, N4910, N637);
not NOT1 (N4915, N4905);
buf BUF1 (N4916, N4908);
not NOT1 (N4917, N4907);
buf BUF1 (N4918, N4901);
or OR4 (N4919, N4912, N4699, N2304, N3831);
or OR4 (N4920, N4911, N3020, N1818, N1014);
and AND4 (N4921, N4914, N3369, N974, N3289);
nor NOR3 (N4922, N4919, N2115, N3573);
xor XOR2 (N4923, N4916, N1426);
buf BUF1 (N4924, N4918);
nor NOR3 (N4925, N4924, N3471, N3128);
nand NAND3 (N4926, N4894, N3041, N2819);
nor NOR3 (N4927, N4917, N4375, N1645);
nor NOR2 (N4928, N4927, N3148);
and AND3 (N4929, N4915, N53, N4905);
not NOT1 (N4930, N4921);
not NOT1 (N4931, N4922);
and AND2 (N4932, N4930, N1589);
xor XOR2 (N4933, N4926, N1090);
xor XOR2 (N4934, N4928, N841);
not NOT1 (N4935, N4923);
xor XOR2 (N4936, N4913, N284);
not NOT1 (N4937, N4920);
nor NOR3 (N4938, N4932, N1316, N2259);
or OR3 (N4939, N4934, N3983, N3671);
or OR4 (N4940, N4903, N4436, N1492, N4264);
or OR2 (N4941, N4936, N826);
not NOT1 (N4942, N4940);
nor NOR2 (N4943, N4941, N338);
or OR2 (N4944, N4937, N170);
buf BUF1 (N4945, N4925);
or OR4 (N4946, N4943, N2692, N1233, N187);
not NOT1 (N4947, N4933);
nand NAND3 (N4948, N4935, N4900, N2015);
xor XOR2 (N4949, N4929, N4103);
not NOT1 (N4950, N4931);
buf BUF1 (N4951, N4947);
xor XOR2 (N4952, N4942, N1336);
xor XOR2 (N4953, N4950, N1815);
or OR3 (N4954, N4939, N3056, N1715);
nor NOR4 (N4955, N4952, N4922, N300, N571);
nor NOR3 (N4956, N4949, N129, N3234);
not NOT1 (N4957, N4956);
buf BUF1 (N4958, N4954);
or OR2 (N4959, N4957, N2182);
xor XOR2 (N4960, N4953, N262);
and AND3 (N4961, N4948, N930, N2119);
or OR2 (N4962, N4955, N2814);
not NOT1 (N4963, N4951);
nor NOR4 (N4964, N4945, N104, N913, N2771);
buf BUF1 (N4965, N4963);
not NOT1 (N4966, N4959);
not NOT1 (N4967, N4964);
not NOT1 (N4968, N4960);
nor NOR3 (N4969, N4968, N4149, N147);
nand NAND3 (N4970, N4938, N1621, N4649);
nor NOR2 (N4971, N4946, N4221);
and AND4 (N4972, N4961, N2664, N2897, N4899);
and AND3 (N4973, N4965, N2951, N4592);
and AND4 (N4974, N4944, N1288, N2166, N2061);
nor NOR2 (N4975, N4962, N479);
nor NOR3 (N4976, N4966, N1385, N1509);
and AND2 (N4977, N4970, N1712);
or OR2 (N4978, N4958, N3246);
or OR4 (N4979, N4971, N561, N4258, N2256);
nand NAND4 (N4980, N4975, N1579, N1798, N789);
nand NAND4 (N4981, N4976, N1680, N1425, N4849);
and AND2 (N4982, N4969, N4696);
xor XOR2 (N4983, N4973, N1126);
buf BUF1 (N4984, N4972);
buf BUF1 (N4985, N4978);
or OR3 (N4986, N4985, N1230, N430);
nand NAND2 (N4987, N4986, N2237);
nand NAND4 (N4988, N4984, N4432, N4851, N2284);
not NOT1 (N4989, N4979);
xor XOR2 (N4990, N4981, N4909);
nor NOR2 (N4991, N4967, N588);
xor XOR2 (N4992, N4983, N2900);
xor XOR2 (N4993, N4980, N4885);
and AND3 (N4994, N4990, N4853, N1091);
nor NOR4 (N4995, N4977, N4675, N3121, N809);
or OR3 (N4996, N4995, N3818, N3505);
not NOT1 (N4997, N4992);
xor XOR2 (N4998, N4974, N1371);
nand NAND3 (N4999, N4988, N631, N1717);
buf BUF1 (N5000, N4999);
nand NAND2 (N5001, N4994, N4842);
nand NAND4 (N5002, N4997, N2162, N4008, N3148);
buf BUF1 (N5003, N4996);
not NOT1 (N5004, N5001);
and AND4 (N5005, N5004, N1922, N966, N4707);
nor NOR3 (N5006, N4991, N2756, N1646);
xor XOR2 (N5007, N4987, N917);
nand NAND2 (N5008, N4993, N198);
nor NOR3 (N5009, N5003, N4356, N1454);
xor XOR2 (N5010, N5002, N13);
or OR2 (N5011, N5005, N4680);
xor XOR2 (N5012, N5010, N4642);
or OR3 (N5013, N4998, N356, N1294);
not NOT1 (N5014, N5009);
and AND2 (N5015, N5008, N3919);
nor NOR4 (N5016, N5015, N1067, N3043, N383);
xor XOR2 (N5017, N4982, N1727);
nand NAND2 (N5018, N5011, N4844);
and AND2 (N5019, N5017, N2032);
nand NAND2 (N5020, N5019, N2814);
nor NOR4 (N5021, N5006, N3131, N4353, N3536);
and AND2 (N5022, N5007, N3156);
or OR3 (N5023, N5013, N1306, N652);
nand NAND3 (N5024, N4989, N2364, N3183);
buf BUF1 (N5025, N5014);
not NOT1 (N5026, N5018);
nand NAND4 (N5027, N5024, N422, N617, N3087);
and AND3 (N5028, N5020, N1863, N1389);
nand NAND3 (N5029, N5028, N1827, N3773);
nand NAND4 (N5030, N5016, N882, N3350, N1803);
not NOT1 (N5031, N5027);
and AND4 (N5032, N5026, N78, N1696, N838);
xor XOR2 (N5033, N5032, N1958);
nor NOR3 (N5034, N5023, N1750, N3422);
and AND4 (N5035, N5031, N3521, N3786, N694);
or OR4 (N5036, N5012, N2541, N191, N1119);
and AND3 (N5037, N5000, N1640, N1888);
not NOT1 (N5038, N5033);
or OR3 (N5039, N5021, N2139, N5016);
not NOT1 (N5040, N5039);
xor XOR2 (N5041, N5034, N1185);
not NOT1 (N5042, N5029);
xor XOR2 (N5043, N5025, N1285);
nand NAND3 (N5044, N5030, N2193, N2449);
nor NOR3 (N5045, N5042, N4033, N4605);
and AND3 (N5046, N5043, N657, N3428);
not NOT1 (N5047, N5046);
nand NAND3 (N5048, N5044, N2985, N4358);
xor XOR2 (N5049, N5035, N3804);
not NOT1 (N5050, N5040);
nor NOR3 (N5051, N5050, N4501, N2542);
not NOT1 (N5052, N5037);
not NOT1 (N5053, N5038);
and AND3 (N5054, N5048, N4550, N3444);
and AND3 (N5055, N5049, N1286, N2905);
and AND2 (N5056, N5045, N4929);
or OR3 (N5057, N5055, N3159, N45);
nand NAND3 (N5058, N5056, N3406, N605);
or OR4 (N5059, N5047, N715, N3258, N613);
or OR2 (N5060, N5052, N941);
xor XOR2 (N5061, N5058, N2583);
or OR2 (N5062, N5059, N347);
not NOT1 (N5063, N5060);
nand NAND4 (N5064, N5036, N1366, N1870, N638);
not NOT1 (N5065, N5064);
or OR2 (N5066, N5065, N648);
buf BUF1 (N5067, N5053);
or OR2 (N5068, N5067, N2371);
xor XOR2 (N5069, N5051, N690);
buf BUF1 (N5070, N5062);
buf BUF1 (N5071, N5063);
or OR3 (N5072, N5070, N1009, N2993);
and AND4 (N5073, N5054, N2791, N4147, N3608);
nand NAND2 (N5074, N5073, N4090);
xor XOR2 (N5075, N5022, N628);
nor NOR4 (N5076, N5041, N2019, N2484, N1284);
nor NOR2 (N5077, N5072, N3132);
or OR4 (N5078, N5069, N1189, N3437, N4078);
buf BUF1 (N5079, N5071);
nor NOR2 (N5080, N5066, N3566);
not NOT1 (N5081, N5061);
not NOT1 (N5082, N5057);
buf BUF1 (N5083, N5078);
buf BUF1 (N5084, N5081);
buf BUF1 (N5085, N5077);
and AND2 (N5086, N5075, N4301);
and AND3 (N5087, N5079, N1009, N1559);
nand NAND2 (N5088, N5084, N2672);
nor NOR2 (N5089, N5085, N1216);
xor XOR2 (N5090, N5087, N19);
not NOT1 (N5091, N5090);
nand NAND2 (N5092, N5080, N2586);
and AND2 (N5093, N5068, N1981);
nor NOR2 (N5094, N5088, N3169);
xor XOR2 (N5095, N5092, N2025);
buf BUF1 (N5096, N5086);
nand NAND4 (N5097, N5095, N4612, N3255, N3913);
and AND3 (N5098, N5091, N2223, N695);
nand NAND4 (N5099, N5098, N226, N830, N2079);
xor XOR2 (N5100, N5097, N3795);
nand NAND2 (N5101, N5082, N550);
and AND2 (N5102, N5096, N3036);
or OR3 (N5103, N5099, N1450, N2749);
xor XOR2 (N5104, N5101, N682);
not NOT1 (N5105, N5093);
and AND4 (N5106, N5104, N2534, N3966, N4967);
or OR2 (N5107, N5094, N2290);
nand NAND4 (N5108, N5103, N2071, N4083, N60);
xor XOR2 (N5109, N5083, N3617);
buf BUF1 (N5110, N5074);
not NOT1 (N5111, N5107);
xor XOR2 (N5112, N5102, N4711);
not NOT1 (N5113, N5076);
not NOT1 (N5114, N5100);
xor XOR2 (N5115, N5105, N2006);
buf BUF1 (N5116, N5110);
not NOT1 (N5117, N5106);
buf BUF1 (N5118, N5113);
nand NAND3 (N5119, N5111, N3270, N2378);
nor NOR2 (N5120, N5115, N4227);
nand NAND4 (N5121, N5089, N2784, N983, N3496);
or OR4 (N5122, N5121, N3381, N3814, N2176);
or OR2 (N5123, N5112, N2439);
or OR2 (N5124, N5122, N341);
xor XOR2 (N5125, N5124, N4964);
and AND3 (N5126, N5116, N1365, N438);
xor XOR2 (N5127, N5119, N2203);
nand NAND4 (N5128, N5108, N3462, N3570, N322);
xor XOR2 (N5129, N5109, N496);
and AND2 (N5130, N5123, N3864);
xor XOR2 (N5131, N5129, N4368);
buf BUF1 (N5132, N5118);
nand NAND4 (N5133, N5125, N1039, N289, N3883);
xor XOR2 (N5134, N5131, N1506);
nor NOR4 (N5135, N5128, N2370, N765, N384);
nand NAND4 (N5136, N5130, N2606, N3730, N4697);
nor NOR2 (N5137, N5135, N1233);
or OR4 (N5138, N5133, N1694, N228, N1244);
buf BUF1 (N5139, N5138);
and AND4 (N5140, N5126, N2369, N1121, N4933);
xor XOR2 (N5141, N5127, N16);
nor NOR4 (N5142, N5114, N2140, N2427, N1385);
or OR4 (N5143, N5136, N4699, N1276, N1994);
buf BUF1 (N5144, N5143);
buf BUF1 (N5145, N5139);
buf BUF1 (N5146, N5134);
nor NOR2 (N5147, N5146, N1105);
nand NAND2 (N5148, N5144, N4546);
nand NAND4 (N5149, N5147, N3540, N2800, N630);
nor NOR4 (N5150, N5132, N4066, N2982, N3364);
buf BUF1 (N5151, N5117);
not NOT1 (N5152, N5151);
xor XOR2 (N5153, N5120, N3761);
nand NAND2 (N5154, N5150, N3927);
or OR4 (N5155, N5153, N4365, N1204, N2093);
not NOT1 (N5156, N5152);
and AND4 (N5157, N5148, N736, N1765, N2618);
and AND3 (N5158, N5140, N3929, N5032);
buf BUF1 (N5159, N5149);
buf BUF1 (N5160, N5142);
and AND4 (N5161, N5137, N3292, N3670, N3050);
nor NOR2 (N5162, N5157, N1703);
nand NAND3 (N5163, N5154, N493, N3214);
or OR3 (N5164, N5163, N1070, N111);
not NOT1 (N5165, N5161);
xor XOR2 (N5166, N5160, N4310);
xor XOR2 (N5167, N5156, N1139);
not NOT1 (N5168, N5165);
xor XOR2 (N5169, N5164, N3179);
and AND2 (N5170, N5162, N3523);
not NOT1 (N5171, N5158);
not NOT1 (N5172, N5141);
and AND2 (N5173, N5155, N1795);
nor NOR3 (N5174, N5170, N2334, N210);
or OR3 (N5175, N5169, N3663, N4764);
xor XOR2 (N5176, N5167, N570);
and AND2 (N5177, N5174, N4235);
nor NOR2 (N5178, N5145, N832);
buf BUF1 (N5179, N5159);
nor NOR2 (N5180, N5175, N3614);
buf BUF1 (N5181, N5176);
xor XOR2 (N5182, N5178, N1313);
nand NAND4 (N5183, N5166, N1561, N5052, N2686);
and AND3 (N5184, N5171, N41, N1126);
and AND3 (N5185, N5168, N3554, N2599);
nor NOR3 (N5186, N5177, N1909, N1995);
buf BUF1 (N5187, N5173);
xor XOR2 (N5188, N5172, N813);
xor XOR2 (N5189, N5188, N3584);
nor NOR2 (N5190, N5187, N1029);
not NOT1 (N5191, N5186);
nand NAND3 (N5192, N5184, N4135, N4688);
and AND3 (N5193, N5180, N3697, N395);
buf BUF1 (N5194, N5182);
and AND2 (N5195, N5194, N1936);
buf BUF1 (N5196, N5195);
buf BUF1 (N5197, N5183);
not NOT1 (N5198, N5197);
not NOT1 (N5199, N5189);
nor NOR2 (N5200, N5181, N2549);
not NOT1 (N5201, N5198);
and AND3 (N5202, N5185, N2191, N1871);
nor NOR3 (N5203, N5193, N1671, N4420);
buf BUF1 (N5204, N5200);
nand NAND2 (N5205, N5190, N1775);
or OR2 (N5206, N5204, N2106);
buf BUF1 (N5207, N5192);
not NOT1 (N5208, N5179);
buf BUF1 (N5209, N5199);
not NOT1 (N5210, N5208);
xor XOR2 (N5211, N5201, N1557);
nor NOR3 (N5212, N5209, N2967, N5152);
buf BUF1 (N5213, N5206);
nor NOR2 (N5214, N5191, N4576);
or OR3 (N5215, N5196, N929, N3211);
or OR2 (N5216, N5211, N3620);
xor XOR2 (N5217, N5205, N52);
xor XOR2 (N5218, N5216, N4340);
buf BUF1 (N5219, N5212);
xor XOR2 (N5220, N5215, N334);
or OR4 (N5221, N5214, N2814, N1560, N2279);
nand NAND3 (N5222, N5202, N3957, N4691);
nor NOR3 (N5223, N5218, N4363, N975);
and AND3 (N5224, N5222, N2269, N2254);
and AND4 (N5225, N5223, N4105, N366, N4392);
xor XOR2 (N5226, N5207, N250);
buf BUF1 (N5227, N5224);
nor NOR2 (N5228, N5226, N4896);
not NOT1 (N5229, N5221);
xor XOR2 (N5230, N5228, N3447);
and AND2 (N5231, N5229, N5091);
buf BUF1 (N5232, N5231);
and AND3 (N5233, N5230, N2878, N1033);
nor NOR4 (N5234, N5225, N984, N2351, N3743);
xor XOR2 (N5235, N5217, N1495);
buf BUF1 (N5236, N5210);
nand NAND3 (N5237, N5236, N148, N1808);
not NOT1 (N5238, N5220);
nand NAND2 (N5239, N5232, N3083);
xor XOR2 (N5240, N5235, N2081);
nor NOR2 (N5241, N5239, N1531);
buf BUF1 (N5242, N5234);
nor NOR4 (N5243, N5237, N539, N1983, N3926);
nor NOR4 (N5244, N5240, N3772, N5192, N2931);
buf BUF1 (N5245, N5227);
nor NOR4 (N5246, N5219, N1789, N3377, N498);
not NOT1 (N5247, N5241);
nor NOR2 (N5248, N5233, N3853);
or OR2 (N5249, N5242, N1831);
buf BUF1 (N5250, N5244);
nand NAND3 (N5251, N5250, N1711, N4650);
nor NOR2 (N5252, N5249, N2801);
not NOT1 (N5253, N5203);
and AND3 (N5254, N5252, N3400, N3715);
and AND4 (N5255, N5253, N1790, N830, N3219);
buf BUF1 (N5256, N5255);
nand NAND4 (N5257, N5243, N4526, N1719, N2027);
nor NOR3 (N5258, N5246, N4930, N4808);
not NOT1 (N5259, N5248);
not NOT1 (N5260, N5251);
nand NAND2 (N5261, N5245, N2657);
buf BUF1 (N5262, N5259);
nor NOR3 (N5263, N5247, N1284, N4733);
or OR2 (N5264, N5260, N4526);
and AND4 (N5265, N5261, N5034, N3685, N3857);
xor XOR2 (N5266, N5262, N2041);
or OR4 (N5267, N5257, N996, N5015, N1320);
and AND2 (N5268, N5213, N1523);
buf BUF1 (N5269, N5268);
not NOT1 (N5270, N5269);
not NOT1 (N5271, N5254);
or OR4 (N5272, N5264, N381, N2940, N3171);
nor NOR2 (N5273, N5271, N85);
and AND4 (N5274, N5258, N2594, N2712, N4558);
or OR3 (N5275, N5263, N1637, N1071);
nand NAND3 (N5276, N5266, N4858, N3316);
xor XOR2 (N5277, N5276, N3398);
buf BUF1 (N5278, N5267);
xor XOR2 (N5279, N5256, N530);
or OR3 (N5280, N5273, N5025, N5259);
xor XOR2 (N5281, N5265, N1860);
nor NOR2 (N5282, N5272, N4848);
buf BUF1 (N5283, N5280);
xor XOR2 (N5284, N5279, N1766);
or OR4 (N5285, N5270, N4479, N3408, N1088);
nand NAND4 (N5286, N5277, N2257, N1671, N1275);
buf BUF1 (N5287, N5282);
nor NOR3 (N5288, N5274, N2522, N1127);
buf BUF1 (N5289, N5284);
or OR3 (N5290, N5275, N3408, N1096);
nand NAND2 (N5291, N5288, N3518);
and AND4 (N5292, N5286, N71, N128, N4607);
not NOT1 (N5293, N5287);
not NOT1 (N5294, N5291);
xor XOR2 (N5295, N5281, N244);
buf BUF1 (N5296, N5294);
buf BUF1 (N5297, N5296);
and AND3 (N5298, N5289, N3311, N3630);
not NOT1 (N5299, N5292);
buf BUF1 (N5300, N5299);
nor NOR4 (N5301, N5283, N2274, N1668, N2873);
xor XOR2 (N5302, N5290, N1300);
and AND4 (N5303, N5301, N2288, N1056, N4059);
xor XOR2 (N5304, N5285, N2185);
nor NOR3 (N5305, N5297, N3364, N2136);
xor XOR2 (N5306, N5298, N559);
or OR2 (N5307, N5305, N4265);
xor XOR2 (N5308, N5293, N3426);
or OR2 (N5309, N5238, N3632);
nand NAND3 (N5310, N5307, N3389, N4391);
nand NAND3 (N5311, N5310, N1015, N577);
buf BUF1 (N5312, N5300);
not NOT1 (N5313, N5278);
xor XOR2 (N5314, N5313, N1239);
and AND2 (N5315, N5306, N3274);
buf BUF1 (N5316, N5309);
or OR3 (N5317, N5304, N895, N2817);
xor XOR2 (N5318, N5303, N2061);
xor XOR2 (N5319, N5302, N1893);
xor XOR2 (N5320, N5314, N837);
xor XOR2 (N5321, N5315, N2798);
nand NAND3 (N5322, N5312, N4872, N2030);
xor XOR2 (N5323, N5321, N1214);
buf BUF1 (N5324, N5311);
nand NAND3 (N5325, N5324, N3484, N4950);
buf BUF1 (N5326, N5316);
or OR2 (N5327, N5317, N4564);
nand NAND4 (N5328, N5326, N4120, N2254, N4851);
or OR3 (N5329, N5295, N2607, N1183);
or OR2 (N5330, N5319, N4901);
and AND2 (N5331, N5322, N3796);
nand NAND3 (N5332, N5308, N885, N5051);
or OR4 (N5333, N5325, N3385, N2398, N4929);
not NOT1 (N5334, N5328);
or OR4 (N5335, N5327, N5271, N1495, N3229);
and AND2 (N5336, N5331, N2986);
xor XOR2 (N5337, N5318, N3489);
nand NAND2 (N5338, N5334, N1610);
nand NAND3 (N5339, N5323, N765, N1893);
xor XOR2 (N5340, N5335, N2510);
or OR2 (N5341, N5330, N4712);
nor NOR2 (N5342, N5341, N3748);
or OR3 (N5343, N5329, N434, N1510);
nand NAND2 (N5344, N5332, N1910);
not NOT1 (N5345, N5340);
nor NOR4 (N5346, N5337, N1533, N1581, N3272);
or OR4 (N5347, N5336, N5293, N2329, N4875);
xor XOR2 (N5348, N5320, N3456);
and AND3 (N5349, N5333, N580, N4399);
xor XOR2 (N5350, N5345, N273);
nor NOR4 (N5351, N5342, N3126, N332, N2591);
nand NAND4 (N5352, N5348, N4666, N5326, N5090);
xor XOR2 (N5353, N5338, N5045);
buf BUF1 (N5354, N5352);
or OR3 (N5355, N5350, N657, N1547);
or OR3 (N5356, N5349, N2648, N2572);
nor NOR3 (N5357, N5346, N2299, N1661);
buf BUF1 (N5358, N5351);
buf BUF1 (N5359, N5344);
and AND3 (N5360, N5356, N4130, N2614);
xor XOR2 (N5361, N5339, N2766);
nand NAND3 (N5362, N5359, N4111, N536);
and AND3 (N5363, N5355, N5112, N3083);
buf BUF1 (N5364, N5347);
buf BUF1 (N5365, N5361);
xor XOR2 (N5366, N5362, N1831);
nor NOR4 (N5367, N5363, N4640, N1006, N737);
not NOT1 (N5368, N5364);
not NOT1 (N5369, N5368);
not NOT1 (N5370, N5354);
xor XOR2 (N5371, N5365, N5370);
or OR3 (N5372, N1961, N4530, N235);
nand NAND4 (N5373, N5372, N5064, N4770, N4958);
not NOT1 (N5374, N5358);
nor NOR3 (N5375, N5367, N5331, N3577);
buf BUF1 (N5376, N5353);
or OR2 (N5377, N5374, N3104);
or OR3 (N5378, N5343, N2276, N849);
or OR4 (N5379, N5375, N2528, N3222, N2998);
and AND2 (N5380, N5366, N4109);
and AND4 (N5381, N5373, N4712, N3545, N1465);
and AND3 (N5382, N5381, N2037, N2356);
not NOT1 (N5383, N5380);
buf BUF1 (N5384, N5360);
or OR4 (N5385, N5383, N3935, N1777, N1159);
nand NAND3 (N5386, N5379, N595, N5003);
xor XOR2 (N5387, N5377, N1234);
and AND2 (N5388, N5376, N293);
and AND4 (N5389, N5371, N5055, N2420, N1477);
buf BUF1 (N5390, N5385);
nand NAND4 (N5391, N5384, N142, N653, N4976);
nand NAND3 (N5392, N5386, N1510, N1578);
nand NAND2 (N5393, N5382, N2336);
or OR3 (N5394, N5389, N3914, N1214);
or OR3 (N5395, N5393, N5356, N4159);
and AND3 (N5396, N5378, N487, N593);
or OR3 (N5397, N5391, N201, N4814);
or OR3 (N5398, N5390, N2222, N1421);
buf BUF1 (N5399, N5395);
buf BUF1 (N5400, N5399);
or OR2 (N5401, N5396, N3771);
buf BUF1 (N5402, N5398);
nor NOR2 (N5403, N5402, N3204);
nand NAND4 (N5404, N5369, N1559, N2782, N3021);
nor NOR4 (N5405, N5388, N3818, N4590, N4242);
nor NOR2 (N5406, N5401, N4663);
or OR2 (N5407, N5405, N1778);
buf BUF1 (N5408, N5406);
nor NOR4 (N5409, N5387, N4854, N2250, N2623);
nor NOR3 (N5410, N5357, N3041, N2378);
nand NAND2 (N5411, N5394, N3981);
or OR4 (N5412, N5408, N5251, N5357, N1347);
not NOT1 (N5413, N5411);
and AND3 (N5414, N5409, N2093, N2617);
not NOT1 (N5415, N5404);
nand NAND2 (N5416, N5413, N4306);
nand NAND4 (N5417, N5403, N3560, N741, N2812);
not NOT1 (N5418, N5407);
or OR2 (N5419, N5412, N3047);
xor XOR2 (N5420, N5416, N1700);
and AND4 (N5421, N5414, N4480, N165, N714);
or OR3 (N5422, N5421, N2804, N2984);
and AND3 (N5423, N5420, N723, N5039);
or OR2 (N5424, N5419, N3100);
or OR2 (N5425, N5400, N2515);
xor XOR2 (N5426, N5422, N773);
and AND3 (N5427, N5417, N1775, N536);
and AND3 (N5428, N5415, N1133, N2667);
nand NAND4 (N5429, N5427, N569, N1791, N3241);
or OR4 (N5430, N5392, N1752, N2726, N1145);
not NOT1 (N5431, N5418);
not NOT1 (N5432, N5397);
nand NAND3 (N5433, N5425, N4798, N2571);
and AND4 (N5434, N5426, N4719, N3226, N2179);
or OR2 (N5435, N5432, N1075);
xor XOR2 (N5436, N5430, N970);
or OR4 (N5437, N5434, N3127, N350, N2958);
xor XOR2 (N5438, N5436, N4149);
nand NAND4 (N5439, N5431, N1495, N3598, N448);
xor XOR2 (N5440, N5424, N4048);
nor NOR2 (N5441, N5440, N2269);
and AND2 (N5442, N5435, N1368);
or OR3 (N5443, N5439, N5067, N1871);
xor XOR2 (N5444, N5441, N4300);
nor NOR4 (N5445, N5442, N4701, N727, N1740);
nor NOR3 (N5446, N5438, N1429, N4518);
nor NOR3 (N5447, N5423, N2429, N5443);
xor XOR2 (N5448, N3422, N2104);
nor NOR2 (N5449, N5445, N4912);
and AND3 (N5450, N5449, N3425, N3420);
nand NAND3 (N5451, N5429, N780, N2022);
not NOT1 (N5452, N5447);
and AND3 (N5453, N5446, N3394, N3233);
nand NAND2 (N5454, N5444, N2912);
or OR4 (N5455, N5428, N864, N5399, N1667);
nor NOR4 (N5456, N5437, N3232, N2569, N1489);
xor XOR2 (N5457, N5455, N2878);
not NOT1 (N5458, N5452);
nor NOR3 (N5459, N5433, N3886, N4935);
or OR3 (N5460, N5410, N1630, N3918);
or OR3 (N5461, N5454, N5065, N4780);
nand NAND2 (N5462, N5450, N1460);
buf BUF1 (N5463, N5461);
or OR2 (N5464, N5457, N2050);
and AND2 (N5465, N5458, N3268);
nor NOR2 (N5466, N5463, N8);
nor NOR2 (N5467, N5459, N3780);
not NOT1 (N5468, N5466);
nor NOR2 (N5469, N5464, N1727);
or OR2 (N5470, N5468, N4008);
nand NAND4 (N5471, N5451, N4584, N2109, N1935);
nand NAND2 (N5472, N5471, N2087);
nand NAND2 (N5473, N5448, N5124);
and AND4 (N5474, N5470, N962, N5209, N98);
xor XOR2 (N5475, N5474, N5144);
nand NAND2 (N5476, N5460, N5227);
xor XOR2 (N5477, N5456, N1759);
or OR4 (N5478, N5469, N4852, N2239, N3444);
and AND3 (N5479, N5462, N495, N4107);
nand NAND2 (N5480, N5476, N4898);
not NOT1 (N5481, N5477);
xor XOR2 (N5482, N5478, N858);
and AND2 (N5483, N5479, N2323);
not NOT1 (N5484, N5482);
and AND2 (N5485, N5481, N2360);
buf BUF1 (N5486, N5465);
xor XOR2 (N5487, N5467, N4240);
buf BUF1 (N5488, N5453);
or OR2 (N5489, N5473, N4644);
and AND3 (N5490, N5489, N519, N4894);
and AND3 (N5491, N5472, N4182, N2849);
buf BUF1 (N5492, N5484);
xor XOR2 (N5493, N5492, N5178);
xor XOR2 (N5494, N5475, N3221);
nor NOR2 (N5495, N5490, N3216);
or OR3 (N5496, N5485, N5078, N2691);
and AND3 (N5497, N5494, N2368, N5246);
nor NOR3 (N5498, N5493, N1363, N4355);
not NOT1 (N5499, N5495);
or OR3 (N5500, N5498, N1072, N1558);
xor XOR2 (N5501, N5480, N5202);
nand NAND3 (N5502, N5499, N330, N3354);
xor XOR2 (N5503, N5486, N3750);
nor NOR4 (N5504, N5483, N2156, N4399, N1595);
and AND2 (N5505, N5504, N5257);
nor NOR2 (N5506, N5487, N4079);
or OR4 (N5507, N5505, N539, N5222, N3814);
not NOT1 (N5508, N5491);
and AND2 (N5509, N5502, N2434);
and AND4 (N5510, N5508, N1070, N86, N3114);
not NOT1 (N5511, N5496);
xor XOR2 (N5512, N5510, N2982);
buf BUF1 (N5513, N5511);
nand NAND2 (N5514, N5507, N3963);
and AND4 (N5515, N5509, N2198, N5358, N882);
buf BUF1 (N5516, N5503);
not NOT1 (N5517, N5516);
not NOT1 (N5518, N5512);
and AND4 (N5519, N5515, N1473, N3143, N1713);
buf BUF1 (N5520, N5513);
or OR2 (N5521, N5497, N2762);
or OR2 (N5522, N5517, N3893);
nor NOR3 (N5523, N5514, N4014, N2089);
or OR4 (N5524, N5500, N559, N5195, N667);
nand NAND4 (N5525, N5501, N432, N927, N4670);
or OR3 (N5526, N5506, N3312, N1099);
xor XOR2 (N5527, N5523, N4145);
xor XOR2 (N5528, N5488, N3323);
xor XOR2 (N5529, N5519, N1558);
and AND4 (N5530, N5529, N2931, N559, N3452);
or OR3 (N5531, N5526, N2680, N46);
not NOT1 (N5532, N5527);
xor XOR2 (N5533, N5530, N1324);
xor XOR2 (N5534, N5528, N683);
xor XOR2 (N5535, N5525, N5430);
not NOT1 (N5536, N5531);
xor XOR2 (N5537, N5524, N838);
nand NAND3 (N5538, N5533, N5183, N1782);
xor XOR2 (N5539, N5520, N852);
and AND2 (N5540, N5518, N5311);
buf BUF1 (N5541, N5540);
nand NAND4 (N5542, N5534, N1988, N478, N2145);
not NOT1 (N5543, N5537);
and AND2 (N5544, N5541, N3892);
xor XOR2 (N5545, N5535, N4927);
not NOT1 (N5546, N5544);
xor XOR2 (N5547, N5521, N3785);
buf BUF1 (N5548, N5542);
nor NOR4 (N5549, N5532, N2370, N1101, N652);
not NOT1 (N5550, N5539);
buf BUF1 (N5551, N5545);
xor XOR2 (N5552, N5550, N2294);
or OR3 (N5553, N5551, N4638, N2876);
and AND4 (N5554, N5543, N25, N4952, N1736);
nand NAND2 (N5555, N5547, N5544);
xor XOR2 (N5556, N5554, N1782);
xor XOR2 (N5557, N5556, N4831);
xor XOR2 (N5558, N5538, N2454);
or OR2 (N5559, N5555, N2180);
not NOT1 (N5560, N5557);
nand NAND2 (N5561, N5548, N970);
not NOT1 (N5562, N5558);
nand NAND4 (N5563, N5536, N1382, N4076, N2065);
and AND2 (N5564, N5549, N4887);
or OR3 (N5565, N5560, N2974, N5507);
not NOT1 (N5566, N5563);
buf BUF1 (N5567, N5522);
buf BUF1 (N5568, N5559);
buf BUF1 (N5569, N5552);
not NOT1 (N5570, N5568);
nor NOR3 (N5571, N5566, N4745, N3380);
xor XOR2 (N5572, N5565, N5244);
xor XOR2 (N5573, N5564, N4875);
or OR2 (N5574, N5567, N1651);
or OR3 (N5575, N5569, N2282, N4541);
xor XOR2 (N5576, N5570, N3506);
or OR2 (N5577, N5561, N3030);
buf BUF1 (N5578, N5546);
nand NAND3 (N5579, N5571, N3344, N1851);
buf BUF1 (N5580, N5575);
or OR4 (N5581, N5576, N726, N775, N369);
nand NAND3 (N5582, N5579, N814, N1339);
xor XOR2 (N5583, N5553, N553);
nand NAND2 (N5584, N5562, N3107);
or OR4 (N5585, N5581, N3918, N5072, N2017);
or OR4 (N5586, N5580, N4773, N2590, N329);
nor NOR2 (N5587, N5578, N449);
not NOT1 (N5588, N5583);
and AND2 (N5589, N5586, N1800);
and AND2 (N5590, N5574, N403);
not NOT1 (N5591, N5584);
or OR2 (N5592, N5585, N5396);
nand NAND4 (N5593, N5592, N3097, N3675, N427);
not NOT1 (N5594, N5587);
xor XOR2 (N5595, N5573, N687);
xor XOR2 (N5596, N5595, N294);
xor XOR2 (N5597, N5594, N2091);
not NOT1 (N5598, N5590);
and AND2 (N5599, N5597, N3697);
buf BUF1 (N5600, N5591);
or OR3 (N5601, N5599, N1846, N1010);
buf BUF1 (N5602, N5588);
not NOT1 (N5603, N5602);
buf BUF1 (N5604, N5603);
nor NOR4 (N5605, N5572, N4738, N612, N2567);
xor XOR2 (N5606, N5605, N3865);
nand NAND3 (N5607, N5577, N1295, N4301);
nand NAND2 (N5608, N5582, N1502);
not NOT1 (N5609, N5604);
nand NAND4 (N5610, N5607, N776, N4349, N2518);
nor NOR4 (N5611, N5609, N4782, N3206, N3282);
buf BUF1 (N5612, N5596);
and AND3 (N5613, N5598, N3801, N5304);
xor XOR2 (N5614, N5606, N1004);
nand NAND3 (N5615, N5612, N5481, N4968);
nor NOR4 (N5616, N5613, N4950, N1971, N3450);
or OR3 (N5617, N5600, N1766, N5516);
nand NAND4 (N5618, N5601, N5005, N3000, N990);
and AND3 (N5619, N5616, N2156, N3519);
and AND4 (N5620, N5615, N2837, N127, N236);
nand NAND2 (N5621, N5614, N2998);
not NOT1 (N5622, N5608);
or OR4 (N5623, N5610, N3721, N4307, N2114);
nor NOR4 (N5624, N5618, N469, N438, N3804);
xor XOR2 (N5625, N5593, N2223);
buf BUF1 (N5626, N5620);
or OR2 (N5627, N5589, N1273);
nor NOR3 (N5628, N5617, N4855, N4916);
or OR4 (N5629, N5627, N4915, N5570, N817);
and AND3 (N5630, N5623, N1709, N3925);
buf BUF1 (N5631, N5629);
or OR2 (N5632, N5630, N1421);
and AND3 (N5633, N5611, N1602, N2944);
buf BUF1 (N5634, N5624);
nor NOR3 (N5635, N5632, N3519, N2333);
and AND2 (N5636, N5622, N953);
nor NOR4 (N5637, N5625, N2036, N1605, N4911);
xor XOR2 (N5638, N5635, N673);
xor XOR2 (N5639, N5628, N4036);
xor XOR2 (N5640, N5621, N3336);
buf BUF1 (N5641, N5638);
or OR2 (N5642, N5634, N1823);
or OR3 (N5643, N5636, N4262, N5183);
not NOT1 (N5644, N5639);
nand NAND3 (N5645, N5643, N4609, N5243);
or OR4 (N5646, N5637, N729, N4650, N2954);
or OR2 (N5647, N5645, N2731);
xor XOR2 (N5648, N5631, N234);
nor NOR2 (N5649, N5619, N2642);
nor NOR3 (N5650, N5648, N427, N3042);
buf BUF1 (N5651, N5649);
xor XOR2 (N5652, N5642, N5377);
and AND2 (N5653, N5640, N5614);
and AND2 (N5654, N5626, N5039);
nand NAND3 (N5655, N5651, N2769, N320);
nand NAND4 (N5656, N5633, N3557, N1858, N495);
and AND4 (N5657, N5644, N5122, N487, N5647);
nand NAND2 (N5658, N2062, N2986);
nand NAND4 (N5659, N5656, N4292, N4531, N2595);
not NOT1 (N5660, N5655);
or OR2 (N5661, N5653, N3385);
nand NAND3 (N5662, N5650, N1605, N140);
nand NAND4 (N5663, N5662, N1761, N4909, N2562);
not NOT1 (N5664, N5663);
nor NOR4 (N5665, N5654, N1121, N5426, N27);
nand NAND2 (N5666, N5660, N1208);
and AND4 (N5667, N5659, N5330, N3743, N488);
and AND2 (N5668, N5664, N1559);
xor XOR2 (N5669, N5665, N2519);
or OR3 (N5670, N5669, N2906, N5382);
or OR2 (N5671, N5657, N4945);
not NOT1 (N5672, N5670);
nand NAND4 (N5673, N5641, N1438, N2254, N2688);
buf BUF1 (N5674, N5668);
buf BUF1 (N5675, N5666);
xor XOR2 (N5676, N5646, N1838);
and AND3 (N5677, N5675, N4094, N3637);
nand NAND4 (N5678, N5652, N956, N1329, N3856);
and AND2 (N5679, N5676, N4220);
or OR3 (N5680, N5671, N2760, N2695);
not NOT1 (N5681, N5678);
nand NAND4 (N5682, N5661, N5204, N4250, N4369);
nand NAND3 (N5683, N5658, N310, N3895);
buf BUF1 (N5684, N5667);
nor NOR4 (N5685, N5683, N33, N4666, N530);
nor NOR2 (N5686, N5674, N1389);
buf BUF1 (N5687, N5677);
xor XOR2 (N5688, N5679, N816);
buf BUF1 (N5689, N5684);
buf BUF1 (N5690, N5689);
nand NAND4 (N5691, N5680, N2415, N2180, N1752);
not NOT1 (N5692, N5685);
not NOT1 (N5693, N5672);
and AND2 (N5694, N5686, N2759);
xor XOR2 (N5695, N5693, N5178);
or OR2 (N5696, N5682, N4806);
nor NOR3 (N5697, N5690, N1492, N5460);
or OR3 (N5698, N5691, N4379, N4558);
nand NAND3 (N5699, N5673, N1439, N3156);
and AND4 (N5700, N5695, N3028, N569, N2652);
and AND2 (N5701, N5688, N5655);
and AND4 (N5702, N5692, N4321, N2600, N2049);
or OR3 (N5703, N5700, N418, N5374);
nor NOR3 (N5704, N5701, N5317, N2800);
and AND3 (N5705, N5697, N4570, N59);
nand NAND3 (N5706, N5699, N3739, N3628);
or OR2 (N5707, N5702, N1709);
buf BUF1 (N5708, N5704);
and AND4 (N5709, N5681, N5308, N5680, N3001);
nand NAND4 (N5710, N5694, N2897, N3703, N2637);
and AND3 (N5711, N5687, N42, N5451);
nand NAND2 (N5712, N5705, N2646);
nor NOR2 (N5713, N5703, N2277);
nor NOR2 (N5714, N5710, N3139);
or OR4 (N5715, N5713, N4112, N3115, N468);
not NOT1 (N5716, N5708);
nand NAND3 (N5717, N5709, N2494, N3301);
and AND4 (N5718, N5714, N4767, N2977, N1919);
not NOT1 (N5719, N5707);
nand NAND2 (N5720, N5717, N5592);
buf BUF1 (N5721, N5698);
nand NAND2 (N5722, N5706, N2070);
xor XOR2 (N5723, N5722, N1130);
buf BUF1 (N5724, N5720);
nand NAND3 (N5725, N5718, N2215, N4743);
or OR2 (N5726, N5725, N5450);
or OR2 (N5727, N5723, N1745);
or OR3 (N5728, N5724, N5287, N4746);
buf BUF1 (N5729, N5719);
nor NOR2 (N5730, N5726, N5670);
buf BUF1 (N5731, N5716);
nor NOR4 (N5732, N5696, N5696, N1068, N1263);
not NOT1 (N5733, N5731);
not NOT1 (N5734, N5711);
nor NOR4 (N5735, N5732, N3150, N226, N1494);
not NOT1 (N5736, N5735);
not NOT1 (N5737, N5727);
nor NOR4 (N5738, N5729, N4979, N3724, N3926);
nand NAND4 (N5739, N5728, N1033, N637, N3886);
xor XOR2 (N5740, N5734, N5379);
nor NOR2 (N5741, N5730, N5599);
and AND2 (N5742, N5738, N5467);
and AND4 (N5743, N5736, N5607, N1644, N3668);
and AND3 (N5744, N5721, N4071, N5339);
nor NOR2 (N5745, N5712, N5621);
and AND2 (N5746, N5741, N955);
nand NAND3 (N5747, N5742, N2818, N3843);
xor XOR2 (N5748, N5733, N443);
xor XOR2 (N5749, N5746, N2164);
or OR4 (N5750, N5747, N3038, N5396, N3422);
or OR2 (N5751, N5743, N3403);
xor XOR2 (N5752, N5748, N4808);
not NOT1 (N5753, N5739);
nor NOR4 (N5754, N5750, N5621, N816, N2442);
xor XOR2 (N5755, N5749, N3208);
and AND4 (N5756, N5754, N5583, N5694, N3325);
not NOT1 (N5757, N5753);
or OR4 (N5758, N5740, N2660, N2983, N3917);
or OR3 (N5759, N5757, N2009, N4184);
not NOT1 (N5760, N5715);
not NOT1 (N5761, N5759);
nor NOR2 (N5762, N5745, N2893);
buf BUF1 (N5763, N5760);
xor XOR2 (N5764, N5756, N3001);
buf BUF1 (N5765, N5752);
buf BUF1 (N5766, N5737);
not NOT1 (N5767, N5764);
not NOT1 (N5768, N5761);
xor XOR2 (N5769, N5758, N3019);
not NOT1 (N5770, N5769);
nand NAND4 (N5771, N5751, N3815, N3526, N4185);
and AND4 (N5772, N5768, N2815, N4950, N868);
or OR2 (N5773, N5744, N4583);
and AND3 (N5774, N5767, N4253, N737);
nand NAND3 (N5775, N5773, N1002, N3248);
nor NOR2 (N5776, N5771, N1316);
buf BUF1 (N5777, N5776);
not NOT1 (N5778, N5774);
or OR2 (N5779, N5762, N2208);
nor NOR4 (N5780, N5778, N3027, N2760, N86);
xor XOR2 (N5781, N5770, N3541);
and AND3 (N5782, N5755, N1087, N3708);
and AND3 (N5783, N5781, N4101, N1841);
not NOT1 (N5784, N5783);
xor XOR2 (N5785, N5766, N4009);
nand NAND3 (N5786, N5785, N1167, N1343);
buf BUF1 (N5787, N5763);
buf BUF1 (N5788, N5787);
and AND4 (N5789, N5788, N69, N5103, N4814);
and AND2 (N5790, N5786, N812);
and AND4 (N5791, N5777, N2267, N1986, N817);
or OR4 (N5792, N5789, N770, N779, N1921);
not NOT1 (N5793, N5791);
and AND2 (N5794, N5775, N2832);
or OR3 (N5795, N5772, N2546, N4960);
buf BUF1 (N5796, N5784);
nor NOR4 (N5797, N5795, N4062, N4073, N4649);
nand NAND3 (N5798, N5794, N2935, N2287);
or OR2 (N5799, N5797, N241);
and AND4 (N5800, N5793, N5457, N4745, N5749);
and AND2 (N5801, N5800, N1405);
not NOT1 (N5802, N5798);
or OR3 (N5803, N5802, N4960, N5007);
and AND4 (N5804, N5801, N4613, N5695, N3836);
nor NOR4 (N5805, N5765, N1844, N2556, N1548);
or OR4 (N5806, N5792, N105, N4047, N1656);
buf BUF1 (N5807, N5805);
or OR3 (N5808, N5806, N1092, N2443);
nor NOR2 (N5809, N5796, N129);
xor XOR2 (N5810, N5804, N3187);
nor NOR3 (N5811, N5810, N706, N3900);
xor XOR2 (N5812, N5809, N1137);
not NOT1 (N5813, N5799);
not NOT1 (N5814, N5780);
xor XOR2 (N5815, N5808, N58);
or OR3 (N5816, N5803, N4613, N5419);
not NOT1 (N5817, N5790);
buf BUF1 (N5818, N5817);
xor XOR2 (N5819, N5813, N2540);
buf BUF1 (N5820, N5779);
nand NAND4 (N5821, N5816, N64, N2775, N4436);
nor NOR3 (N5822, N5782, N5557, N830);
not NOT1 (N5823, N5807);
and AND4 (N5824, N5822, N4080, N3783, N83);
and AND3 (N5825, N5811, N3023, N1326);
xor XOR2 (N5826, N5818, N4343);
or OR4 (N5827, N5819, N5748, N4500, N1571);
nor NOR4 (N5828, N5815, N1757, N2661, N856);
or OR4 (N5829, N5820, N4209, N3271, N3340);
buf BUF1 (N5830, N5826);
not NOT1 (N5831, N5828);
and AND2 (N5832, N5830, N5776);
xor XOR2 (N5833, N5832, N5122);
not NOT1 (N5834, N5825);
or OR3 (N5835, N5827, N863, N99);
xor XOR2 (N5836, N5824, N2212);
nand NAND3 (N5837, N5829, N2154, N1678);
xor XOR2 (N5838, N5823, N4652);
or OR2 (N5839, N5835, N1099);
buf BUF1 (N5840, N5839);
not NOT1 (N5841, N5840);
nor NOR4 (N5842, N5836, N5714, N898, N1185);
not NOT1 (N5843, N5833);
xor XOR2 (N5844, N5834, N4314);
not NOT1 (N5845, N5831);
and AND4 (N5846, N5843, N1611, N2320, N5701);
nor NOR3 (N5847, N5821, N770, N1103);
nor NOR2 (N5848, N5847, N680);
not NOT1 (N5849, N5812);
not NOT1 (N5850, N5842);
nand NAND2 (N5851, N5844, N1135);
or OR3 (N5852, N5851, N2285, N107);
not NOT1 (N5853, N5852);
nand NAND3 (N5854, N5841, N1422, N2284);
nand NAND3 (N5855, N5837, N993, N1578);
and AND2 (N5856, N5855, N3050);
not NOT1 (N5857, N5849);
xor XOR2 (N5858, N5845, N1546);
nor NOR4 (N5859, N5814, N4630, N609, N1584);
not NOT1 (N5860, N5850);
nand NAND3 (N5861, N5856, N636, N4412);
not NOT1 (N5862, N5859);
buf BUF1 (N5863, N5853);
buf BUF1 (N5864, N5860);
nand NAND3 (N5865, N5854, N5363, N1605);
xor XOR2 (N5866, N5862, N4415);
not NOT1 (N5867, N5846);
not NOT1 (N5868, N5848);
and AND3 (N5869, N5867, N4797, N1825);
not NOT1 (N5870, N5864);
nor NOR4 (N5871, N5868, N3682, N1270, N4603);
not NOT1 (N5872, N5863);
and AND3 (N5873, N5838, N2359, N3872);
nand NAND3 (N5874, N5866, N4579, N2486);
not NOT1 (N5875, N5865);
nand NAND4 (N5876, N5872, N1322, N655, N1890);
and AND2 (N5877, N5875, N3225);
nor NOR4 (N5878, N5877, N3827, N2134, N112);
buf BUF1 (N5879, N5861);
nand NAND3 (N5880, N5857, N3714, N4181);
nand NAND2 (N5881, N5879, N5302);
and AND2 (N5882, N5881, N3023);
xor XOR2 (N5883, N5880, N2672);
and AND2 (N5884, N5873, N4683);
buf BUF1 (N5885, N5858);
xor XOR2 (N5886, N5876, N5145);
not NOT1 (N5887, N5885);
or OR2 (N5888, N5869, N3597);
xor XOR2 (N5889, N5874, N4437);
nand NAND2 (N5890, N5870, N4492);
xor XOR2 (N5891, N5890, N4579);
xor XOR2 (N5892, N5883, N2387);
buf BUF1 (N5893, N5882);
xor XOR2 (N5894, N5887, N4688);
xor XOR2 (N5895, N5894, N4577);
and AND4 (N5896, N5878, N1429, N3075, N925);
nor NOR4 (N5897, N5884, N4268, N1859, N2170);
not NOT1 (N5898, N5871);
and AND4 (N5899, N5893, N5127, N1900, N2696);
not NOT1 (N5900, N5897);
and AND4 (N5901, N5888, N3419, N3426, N4155);
or OR2 (N5902, N5895, N1314);
or OR4 (N5903, N5896, N2603, N4820, N5531);
nor NOR3 (N5904, N5901, N655, N48);
not NOT1 (N5905, N5898);
not NOT1 (N5906, N5892);
or OR4 (N5907, N5900, N4651, N5576, N3089);
and AND3 (N5908, N5907, N291, N494);
nand NAND4 (N5909, N5906, N3460, N2269, N4642);
or OR4 (N5910, N5891, N2510, N2262, N3048);
or OR4 (N5911, N5909, N5006, N154, N885);
not NOT1 (N5912, N5902);
nand NAND3 (N5913, N5886, N425, N4339);
or OR2 (N5914, N5905, N1697);
or OR4 (N5915, N5903, N5101, N4150, N4561);
buf BUF1 (N5916, N5915);
or OR3 (N5917, N5914, N3192, N651);
or OR2 (N5918, N5911, N5872);
xor XOR2 (N5919, N5912, N820);
nor NOR2 (N5920, N5913, N3681);
nand NAND3 (N5921, N5918, N4370, N3512);
buf BUF1 (N5922, N5904);
not NOT1 (N5923, N5908);
nor NOR2 (N5924, N5923, N2855);
buf BUF1 (N5925, N5919);
and AND2 (N5926, N5925, N2923);
or OR2 (N5927, N5917, N3900);
nor NOR2 (N5928, N5920, N692);
xor XOR2 (N5929, N5928, N4371);
nand NAND2 (N5930, N5922, N845);
nor NOR2 (N5931, N5910, N4438);
not NOT1 (N5932, N5916);
xor XOR2 (N5933, N5927, N3609);
nand NAND4 (N5934, N5924, N150, N3991, N767);
nor NOR3 (N5935, N5926, N3279, N4903);
not NOT1 (N5936, N5932);
and AND4 (N5937, N5889, N977, N5601, N5373);
nand NAND4 (N5938, N5930, N1872, N5431, N4283);
xor XOR2 (N5939, N5938, N5540);
nand NAND2 (N5940, N5934, N2777);
buf BUF1 (N5941, N5933);
and AND2 (N5942, N5936, N4508);
not NOT1 (N5943, N5935);
and AND3 (N5944, N5940, N4991, N1824);
buf BUF1 (N5945, N5943);
buf BUF1 (N5946, N5945);
buf BUF1 (N5947, N5946);
nand NAND4 (N5948, N5941, N2940, N5229, N1929);
nand NAND4 (N5949, N5947, N2188, N4946, N4686);
not NOT1 (N5950, N5948);
not NOT1 (N5951, N5921);
buf BUF1 (N5952, N5950);
xor XOR2 (N5953, N5939, N1473);
and AND2 (N5954, N5937, N239);
or OR2 (N5955, N5952, N4852);
nor NOR4 (N5956, N5931, N3632, N5909, N1982);
buf BUF1 (N5957, N5949);
nand NAND4 (N5958, N5942, N2641, N1790, N2864);
buf BUF1 (N5959, N5955);
buf BUF1 (N5960, N5956);
not NOT1 (N5961, N5958);
buf BUF1 (N5962, N5929);
buf BUF1 (N5963, N5960);
nand NAND2 (N5964, N5951, N5765);
or OR3 (N5965, N5953, N1739, N4246);
not NOT1 (N5966, N5959);
or OR4 (N5967, N5966, N206, N16, N5335);
nor NOR3 (N5968, N5965, N5661, N5258);
buf BUF1 (N5969, N5961);
nand NAND2 (N5970, N5968, N2678);
or OR2 (N5971, N5967, N1549);
nand NAND2 (N5972, N5944, N3056);
nor NOR4 (N5973, N5963, N2131, N1634, N20);
or OR2 (N5974, N5970, N2667);
or OR2 (N5975, N5973, N1088);
and AND3 (N5976, N5971, N2055, N5966);
nand NAND3 (N5977, N5954, N5941, N1913);
and AND4 (N5978, N5976, N5080, N4086, N1221);
nand NAND4 (N5979, N5978, N2808, N676, N910);
or OR2 (N5980, N5899, N5194);
not NOT1 (N5981, N5980);
not NOT1 (N5982, N5969);
buf BUF1 (N5983, N5972);
not NOT1 (N5984, N5957);
and AND3 (N5985, N5975, N2028, N4505);
not NOT1 (N5986, N5962);
buf BUF1 (N5987, N5979);
nand NAND3 (N5988, N5974, N3749, N3929);
and AND3 (N5989, N5983, N1690, N801);
and AND3 (N5990, N5988, N4572, N5173);
not NOT1 (N5991, N5985);
or OR3 (N5992, N5991, N3537, N2459);
or OR3 (N5993, N5964, N109, N3964);
not NOT1 (N5994, N5989);
xor XOR2 (N5995, N5990, N3016);
xor XOR2 (N5996, N5977, N3906);
nor NOR4 (N5997, N5994, N4428, N5241, N995);
xor XOR2 (N5998, N5997, N544);
not NOT1 (N5999, N5981);
not NOT1 (N6000, N5986);
or OR2 (N6001, N6000, N4821);
buf BUF1 (N6002, N5993);
nor NOR3 (N6003, N5982, N5990, N2432);
nand NAND3 (N6004, N5998, N3137, N221);
xor XOR2 (N6005, N5984, N1926);
buf BUF1 (N6006, N5999);
buf BUF1 (N6007, N6001);
and AND3 (N6008, N5995, N3230, N1482);
or OR2 (N6009, N6004, N4444);
or OR3 (N6010, N6005, N3145, N332);
not NOT1 (N6011, N6003);
buf BUF1 (N6012, N5987);
or OR4 (N6013, N6002, N561, N940, N5392);
not NOT1 (N6014, N6008);
or OR2 (N6015, N6010, N2836);
xor XOR2 (N6016, N6011, N5888);
not NOT1 (N6017, N6009);
nand NAND2 (N6018, N5992, N2164);
buf BUF1 (N6019, N5996);
and AND3 (N6020, N6012, N1303, N4784);
xor XOR2 (N6021, N6018, N21);
nor NOR2 (N6022, N6017, N4284);
xor XOR2 (N6023, N6013, N4521);
not NOT1 (N6024, N6020);
xor XOR2 (N6025, N6023, N5649);
and AND3 (N6026, N6006, N3224, N2809);
xor XOR2 (N6027, N6025, N985);
buf BUF1 (N6028, N6007);
nor NOR2 (N6029, N6015, N934);
nor NOR3 (N6030, N6028, N2126, N146);
and AND2 (N6031, N6014, N5363);
buf BUF1 (N6032, N6016);
not NOT1 (N6033, N6029);
and AND3 (N6034, N6024, N3211, N5244);
nor NOR3 (N6035, N6032, N473, N5598);
not NOT1 (N6036, N6035);
and AND2 (N6037, N6030, N1825);
and AND4 (N6038, N6026, N1974, N855, N4054);
xor XOR2 (N6039, N6022, N1009);
or OR2 (N6040, N6038, N4421);
nor NOR3 (N6041, N6039, N5325, N2047);
nor NOR2 (N6042, N6040, N2448);
nor NOR4 (N6043, N6036, N1722, N3901, N1418);
nor NOR4 (N6044, N6021, N4908, N4318, N4404);
nor NOR3 (N6045, N6043, N2024, N2401);
xor XOR2 (N6046, N6042, N2521);
nor NOR2 (N6047, N6044, N3057);
nand NAND2 (N6048, N6047, N1412);
and AND3 (N6049, N6033, N477, N5546);
not NOT1 (N6050, N6037);
nand NAND3 (N6051, N6048, N3469, N6007);
and AND2 (N6052, N6049, N451);
not NOT1 (N6053, N6031);
and AND4 (N6054, N6046, N1169, N5590, N2657);
nor NOR4 (N6055, N6045, N3628, N1229, N25);
buf BUF1 (N6056, N6019);
xor XOR2 (N6057, N6054, N5081);
or OR4 (N6058, N6051, N5986, N3122, N4479);
buf BUF1 (N6059, N6053);
nand NAND4 (N6060, N6056, N746, N2168, N1866);
buf BUF1 (N6061, N6059);
buf BUF1 (N6062, N6058);
or OR4 (N6063, N6052, N1225, N5729, N5718);
nor NOR4 (N6064, N6027, N5645, N3413, N2967);
not NOT1 (N6065, N6050);
not NOT1 (N6066, N6063);
nor NOR2 (N6067, N6060, N213);
nand NAND3 (N6068, N6065, N3744, N5395);
nand NAND2 (N6069, N6041, N1232);
and AND4 (N6070, N6062, N1539, N4723, N1987);
or OR2 (N6071, N6070, N1479);
xor XOR2 (N6072, N6066, N3498);
xor XOR2 (N6073, N6069, N1941);
nor NOR3 (N6074, N6073, N5144, N3666);
and AND4 (N6075, N6071, N2171, N3765, N4577);
xor XOR2 (N6076, N6074, N1687);
xor XOR2 (N6077, N6055, N642);
nand NAND4 (N6078, N6057, N1264, N2801, N437);
or OR3 (N6079, N6061, N979, N446);
buf BUF1 (N6080, N6068);
or OR3 (N6081, N6064, N124, N5670);
xor XOR2 (N6082, N6078, N4119);
not NOT1 (N6083, N6080);
xor XOR2 (N6084, N6083, N634);
or OR2 (N6085, N6084, N646);
buf BUF1 (N6086, N6076);
nor NOR4 (N6087, N6085, N4639, N4492, N5046);
buf BUF1 (N6088, N6072);
xor XOR2 (N6089, N6088, N1012);
nand NAND4 (N6090, N6075, N3283, N1164, N1953);
buf BUF1 (N6091, N6067);
nor NOR2 (N6092, N6086, N910);
not NOT1 (N6093, N6090);
nand NAND2 (N6094, N6087, N5130);
buf BUF1 (N6095, N6081);
and AND2 (N6096, N6077, N3687);
buf BUF1 (N6097, N6093);
nand NAND4 (N6098, N6092, N1559, N4087, N1011);
not NOT1 (N6099, N6098);
not NOT1 (N6100, N6095);
nand NAND3 (N6101, N6099, N1249, N3866);
and AND2 (N6102, N6101, N4174);
and AND4 (N6103, N6100, N62, N4926, N2471);
buf BUF1 (N6104, N6094);
xor XOR2 (N6105, N6034, N31);
not NOT1 (N6106, N6082);
nand NAND4 (N6107, N6106, N683, N3378, N4712);
not NOT1 (N6108, N6103);
nand NAND2 (N6109, N6105, N4994);
nor NOR2 (N6110, N6107, N1043);
nand NAND2 (N6111, N6108, N5885);
or OR4 (N6112, N6110, N5069, N1551, N1965);
buf BUF1 (N6113, N6079);
not NOT1 (N6114, N6096);
or OR4 (N6115, N6104, N422, N5599, N4980);
xor XOR2 (N6116, N6111, N5151);
or OR3 (N6117, N6109, N109, N1452);
buf BUF1 (N6118, N6102);
nand NAND3 (N6119, N6113, N1864, N1302);
or OR4 (N6120, N6118, N1779, N1143, N559);
and AND4 (N6121, N6117, N59, N2414, N2496);
xor XOR2 (N6122, N6114, N4138);
nor NOR4 (N6123, N6116, N2152, N901, N562);
nand NAND2 (N6124, N6091, N2697);
buf BUF1 (N6125, N6123);
nor NOR4 (N6126, N6122, N4948, N1764, N3604);
not NOT1 (N6127, N6126);
or OR2 (N6128, N6125, N3568);
nand NAND4 (N6129, N6127, N3063, N3264, N4877);
not NOT1 (N6130, N6115);
nor NOR4 (N6131, N6124, N4209, N1055, N3603);
nand NAND4 (N6132, N6131, N3366, N571, N5844);
and AND4 (N6133, N6128, N3757, N917, N5187);
buf BUF1 (N6134, N6112);
xor XOR2 (N6135, N6132, N3154);
or OR2 (N6136, N6121, N3488);
xor XOR2 (N6137, N6133, N5384);
xor XOR2 (N6138, N6134, N3688);
not NOT1 (N6139, N6135);
nor NOR2 (N6140, N6139, N4125);
not NOT1 (N6141, N6140);
buf BUF1 (N6142, N6129);
and AND4 (N6143, N6137, N3447, N1802, N3570);
not NOT1 (N6144, N6119);
buf BUF1 (N6145, N6144);
and AND3 (N6146, N6097, N2631, N1678);
not NOT1 (N6147, N6089);
buf BUF1 (N6148, N6143);
and AND3 (N6149, N6142, N874, N3209);
and AND2 (N6150, N6145, N2599);
buf BUF1 (N6151, N6150);
nand NAND4 (N6152, N6148, N3490, N544, N397);
buf BUF1 (N6153, N6141);
and AND3 (N6154, N6147, N3845, N92);
nor NOR4 (N6155, N6152, N4039, N6116, N423);
not NOT1 (N6156, N6146);
not NOT1 (N6157, N6153);
and AND3 (N6158, N6154, N4297, N2499);
or OR2 (N6159, N6136, N970);
xor XOR2 (N6160, N6156, N5349);
and AND2 (N6161, N6149, N3340);
nor NOR2 (N6162, N6130, N6);
nor NOR4 (N6163, N6151, N1287, N3805, N5280);
not NOT1 (N6164, N6120);
nand NAND2 (N6165, N6161, N5617);
and AND4 (N6166, N6164, N1363, N1338, N1358);
nor NOR2 (N6167, N6157, N2932);
and AND3 (N6168, N6160, N2463, N3672);
and AND3 (N6169, N6165, N4944, N1043);
not NOT1 (N6170, N6168);
xor XOR2 (N6171, N6170, N1129);
and AND3 (N6172, N6163, N4429, N4525);
not NOT1 (N6173, N6138);
not NOT1 (N6174, N6162);
and AND2 (N6175, N6171, N1007);
and AND3 (N6176, N6175, N6118, N4423);
or OR2 (N6177, N6173, N4617);
buf BUF1 (N6178, N6172);
xor XOR2 (N6179, N6159, N5252);
xor XOR2 (N6180, N6178, N3912);
not NOT1 (N6181, N6155);
and AND4 (N6182, N6169, N788, N3399, N4664);
and AND3 (N6183, N6182, N5457, N3276);
not NOT1 (N6184, N6176);
and AND3 (N6185, N6179, N911, N1388);
nand NAND3 (N6186, N6183, N4795, N3306);
xor XOR2 (N6187, N6158, N6149);
buf BUF1 (N6188, N6174);
buf BUF1 (N6189, N6167);
not NOT1 (N6190, N6185);
nor NOR3 (N6191, N6181, N5982, N5923);
nor NOR3 (N6192, N6166, N3016, N6043);
nor NOR4 (N6193, N6188, N329, N2198, N795);
xor XOR2 (N6194, N6193, N3658);
nor NOR4 (N6195, N6184, N5628, N5025, N4942);
buf BUF1 (N6196, N6177);
xor XOR2 (N6197, N6190, N2113);
nand NAND2 (N6198, N6191, N3729);
not NOT1 (N6199, N6186);
not NOT1 (N6200, N6197);
nand NAND4 (N6201, N6189, N2267, N5660, N70);
and AND2 (N6202, N6194, N5684);
buf BUF1 (N6203, N6198);
and AND3 (N6204, N6201, N873, N2121);
xor XOR2 (N6205, N6187, N5911);
nor NOR2 (N6206, N6203, N3764);
and AND4 (N6207, N6192, N1808, N4381, N3523);
xor XOR2 (N6208, N6207, N2328);
xor XOR2 (N6209, N6208, N5391);
nor NOR4 (N6210, N6200, N1170, N5052, N3021);
and AND3 (N6211, N6180, N3881, N3092);
xor XOR2 (N6212, N6206, N3343);
nor NOR4 (N6213, N6205, N3576, N1500, N1734);
xor XOR2 (N6214, N6204, N1891);
xor XOR2 (N6215, N6199, N5084);
not NOT1 (N6216, N6215);
or OR3 (N6217, N6209, N2676, N5440);
xor XOR2 (N6218, N6214, N5121);
not NOT1 (N6219, N6211);
nor NOR2 (N6220, N6210, N4634);
buf BUF1 (N6221, N6196);
xor XOR2 (N6222, N6213, N455);
and AND2 (N6223, N6220, N2154);
xor XOR2 (N6224, N6218, N2621);
and AND2 (N6225, N6212, N3050);
nand NAND2 (N6226, N6202, N4878);
xor XOR2 (N6227, N6221, N197);
not NOT1 (N6228, N6222);
not NOT1 (N6229, N6225);
xor XOR2 (N6230, N6227, N2474);
nor NOR3 (N6231, N6217, N3983, N2319);
not NOT1 (N6232, N6230);
or OR3 (N6233, N6231, N1763, N3403);
buf BUF1 (N6234, N6224);
not NOT1 (N6235, N6229);
or OR2 (N6236, N6216, N1007);
not NOT1 (N6237, N6232);
xor XOR2 (N6238, N6223, N4007);
or OR4 (N6239, N6228, N1775, N3565, N4055);
not NOT1 (N6240, N6195);
and AND3 (N6241, N6226, N4468, N5525);
and AND4 (N6242, N6219, N1042, N2064, N3518);
nand NAND3 (N6243, N6240, N2651, N37);
or OR2 (N6244, N6243, N5248);
or OR2 (N6245, N6234, N174);
xor XOR2 (N6246, N6241, N1437);
nor NOR3 (N6247, N6236, N3843, N2562);
and AND3 (N6248, N6247, N2513, N1402);
buf BUF1 (N6249, N6245);
nor NOR2 (N6250, N6249, N3361);
buf BUF1 (N6251, N6244);
xor XOR2 (N6252, N6242, N6045);
xor XOR2 (N6253, N6233, N4274);
or OR2 (N6254, N6250, N5065);
and AND2 (N6255, N6238, N811);
or OR2 (N6256, N6255, N6049);
or OR4 (N6257, N6248, N125, N3896, N1242);
xor XOR2 (N6258, N6235, N1088);
or OR2 (N6259, N6251, N940);
buf BUF1 (N6260, N6253);
nor NOR3 (N6261, N6260, N4570, N3897);
xor XOR2 (N6262, N6237, N524);
or OR3 (N6263, N6257, N5570, N341);
xor XOR2 (N6264, N6254, N2471);
xor XOR2 (N6265, N6258, N1936);
nor NOR2 (N6266, N6264, N3749);
buf BUF1 (N6267, N6261);
nand NAND2 (N6268, N6239, N244);
nand NAND2 (N6269, N6267, N5154);
nand NAND3 (N6270, N6268, N808, N6068);
or OR2 (N6271, N6252, N3425);
or OR3 (N6272, N6246, N4322, N2825);
xor XOR2 (N6273, N6271, N945);
xor XOR2 (N6274, N6269, N5674);
and AND4 (N6275, N6272, N2543, N1137, N5701);
not NOT1 (N6276, N6273);
and AND2 (N6277, N6270, N63);
nand NAND3 (N6278, N6256, N752, N2039);
or OR2 (N6279, N6274, N4819);
nand NAND2 (N6280, N6277, N4784);
not NOT1 (N6281, N6276);
buf BUF1 (N6282, N6280);
and AND3 (N6283, N6259, N2749, N4031);
or OR3 (N6284, N6283, N1893, N3023);
or OR2 (N6285, N6284, N4999);
nor NOR4 (N6286, N6278, N1619, N1077, N1821);
buf BUF1 (N6287, N6266);
not NOT1 (N6288, N6287);
or OR3 (N6289, N6275, N134, N4960);
buf BUF1 (N6290, N6281);
and AND2 (N6291, N6282, N465);
not NOT1 (N6292, N6288);
nand NAND4 (N6293, N6265, N949, N5575, N1739);
not NOT1 (N6294, N6291);
buf BUF1 (N6295, N6292);
nor NOR4 (N6296, N6285, N5995, N4777, N1466);
and AND3 (N6297, N6289, N5235, N3910);
nor NOR2 (N6298, N6263, N649);
buf BUF1 (N6299, N6296);
and AND4 (N6300, N6293, N5472, N1073, N2205);
nand NAND3 (N6301, N6297, N5480, N1177);
nor NOR2 (N6302, N6299, N1977);
xor XOR2 (N6303, N6300, N4591);
nand NAND2 (N6304, N6295, N4711);
nor NOR2 (N6305, N6304, N1870);
xor XOR2 (N6306, N6262, N2741);
xor XOR2 (N6307, N6286, N5668);
or OR3 (N6308, N6294, N1361, N2267);
xor XOR2 (N6309, N6302, N5048);
nor NOR3 (N6310, N6309, N611, N5626);
and AND3 (N6311, N6279, N2524, N4745);
or OR3 (N6312, N6311, N2487, N380);
and AND4 (N6313, N6307, N690, N2637, N1956);
nor NOR3 (N6314, N6310, N917, N1996);
xor XOR2 (N6315, N6306, N2477);
or OR2 (N6316, N6305, N4526);
buf BUF1 (N6317, N6301);
and AND2 (N6318, N6315, N3662);
buf BUF1 (N6319, N6316);
not NOT1 (N6320, N6308);
nand NAND4 (N6321, N6318, N1543, N6110, N3634);
buf BUF1 (N6322, N6313);
buf BUF1 (N6323, N6322);
buf BUF1 (N6324, N6312);
or OR4 (N6325, N6319, N594, N2121, N44);
or OR3 (N6326, N6323, N1160, N5524);
not NOT1 (N6327, N6290);
nand NAND2 (N6328, N6298, N521);
not NOT1 (N6329, N6314);
buf BUF1 (N6330, N6320);
nor NOR3 (N6331, N6303, N5940, N150);
xor XOR2 (N6332, N6326, N1613);
or OR3 (N6333, N6324, N922, N5337);
xor XOR2 (N6334, N6329, N3184);
or OR3 (N6335, N6334, N2538, N5073);
nor NOR3 (N6336, N6333, N3835, N752);
and AND3 (N6337, N6335, N4654, N1476);
nor NOR2 (N6338, N6337, N2978);
and AND3 (N6339, N6317, N3647, N1106);
xor XOR2 (N6340, N6325, N5429);
buf BUF1 (N6341, N6336);
nor NOR3 (N6342, N6330, N1335, N2906);
and AND4 (N6343, N6327, N3794, N2968, N4061);
and AND3 (N6344, N6341, N986, N260);
and AND3 (N6345, N6340, N369, N4741);
or OR4 (N6346, N6338, N2047, N881, N5413);
or OR2 (N6347, N6342, N1504);
or OR2 (N6348, N6345, N614);
or OR3 (N6349, N6347, N4875, N5376);
nand NAND3 (N6350, N6346, N3710, N4155);
buf BUF1 (N6351, N6331);
not NOT1 (N6352, N6349);
not NOT1 (N6353, N6332);
nand NAND2 (N6354, N6343, N4769);
or OR4 (N6355, N6348, N3237, N2812, N801);
buf BUF1 (N6356, N6352);
buf BUF1 (N6357, N6350);
and AND3 (N6358, N6353, N1695, N2796);
buf BUF1 (N6359, N6351);
nand NAND2 (N6360, N6359, N322);
buf BUF1 (N6361, N6356);
or OR3 (N6362, N6328, N3828, N3642);
nand NAND2 (N6363, N6355, N1699);
not NOT1 (N6364, N6358);
and AND3 (N6365, N6361, N2930, N3799);
and AND4 (N6366, N6344, N3412, N4042, N1637);
not NOT1 (N6367, N6339);
buf BUF1 (N6368, N6360);
nand NAND4 (N6369, N6368, N5661, N3155, N3036);
not NOT1 (N6370, N6367);
or OR4 (N6371, N6321, N2429, N3301, N386);
nand NAND3 (N6372, N6370, N5096, N3754);
nand NAND2 (N6373, N6357, N4403);
not NOT1 (N6374, N6354);
xor XOR2 (N6375, N6369, N2140);
nor NOR4 (N6376, N6375, N5132, N4508, N1327);
not NOT1 (N6377, N6376);
nand NAND2 (N6378, N6365, N1153);
not NOT1 (N6379, N6378);
and AND4 (N6380, N6364, N3517, N4691, N609);
and AND2 (N6381, N6373, N1141);
nor NOR4 (N6382, N6374, N1294, N4343, N5473);
nor NOR3 (N6383, N6380, N1300, N2690);
and AND2 (N6384, N6372, N4820);
buf BUF1 (N6385, N6362);
xor XOR2 (N6386, N6385, N5508);
nor NOR4 (N6387, N6366, N5406, N4857, N5859);
not NOT1 (N6388, N6377);
or OR3 (N6389, N6382, N2600, N1533);
nor NOR3 (N6390, N6384, N6215, N3753);
or OR4 (N6391, N6390, N3542, N1266, N4104);
xor XOR2 (N6392, N6383, N5154);
xor XOR2 (N6393, N6389, N6197);
or OR2 (N6394, N6391, N5398);
nor NOR3 (N6395, N6387, N119, N1915);
nor NOR2 (N6396, N6381, N811);
nor NOR4 (N6397, N6393, N2048, N2805, N760);
buf BUF1 (N6398, N6396);
nor NOR2 (N6399, N6392, N349);
buf BUF1 (N6400, N6363);
nand NAND3 (N6401, N6398, N2106, N5887);
nor NOR3 (N6402, N6400, N4530, N5098);
not NOT1 (N6403, N6395);
and AND4 (N6404, N6394, N2442, N5700, N3764);
nor NOR3 (N6405, N6399, N1167, N3418);
buf BUF1 (N6406, N6379);
and AND2 (N6407, N6371, N572);
xor XOR2 (N6408, N6388, N987);
buf BUF1 (N6409, N6397);
nor NOR4 (N6410, N6406, N3927, N3472, N3552);
or OR3 (N6411, N6401, N3158, N5260);
nand NAND2 (N6412, N6404, N1365);
nand NAND4 (N6413, N6410, N2251, N5296, N1347);
buf BUF1 (N6414, N6412);
nand NAND3 (N6415, N6403, N118, N4515);
nand NAND2 (N6416, N6413, N5461);
and AND2 (N6417, N6402, N4510);
nand NAND4 (N6418, N6415, N1875, N1451, N2062);
and AND2 (N6419, N6416, N3266);
and AND2 (N6420, N6414, N3375);
nand NAND3 (N6421, N6386, N85, N1771);
nand NAND3 (N6422, N6407, N4253, N3958);
and AND2 (N6423, N6408, N5786);
buf BUF1 (N6424, N6417);
not NOT1 (N6425, N6420);
xor XOR2 (N6426, N6419, N305);
not NOT1 (N6427, N6421);
and AND2 (N6428, N6424, N1309);
buf BUF1 (N6429, N6409);
or OR3 (N6430, N6428, N2869, N4259);
or OR4 (N6431, N6425, N74, N5140, N3690);
nand NAND4 (N6432, N6411, N5321, N5347, N267);
nor NOR2 (N6433, N6423, N3682);
nor NOR2 (N6434, N6429, N1430);
not NOT1 (N6435, N6434);
not NOT1 (N6436, N6435);
not NOT1 (N6437, N6426);
nand NAND4 (N6438, N6437, N3127, N5360, N1419);
not NOT1 (N6439, N6418);
nand NAND3 (N6440, N6427, N1445, N1129);
and AND4 (N6441, N6438, N814, N4392, N2774);
and AND2 (N6442, N6439, N4738);
nor NOR2 (N6443, N6441, N6338);
or OR4 (N6444, N6443, N4685, N3652, N2814);
xor XOR2 (N6445, N6433, N5304);
or OR3 (N6446, N6442, N349, N6317);
xor XOR2 (N6447, N6431, N3609);
or OR2 (N6448, N6432, N4901);
and AND2 (N6449, N6446, N3759);
nor NOR2 (N6450, N6444, N2931);
xor XOR2 (N6451, N6445, N3746);
buf BUF1 (N6452, N6448);
and AND4 (N6453, N6450, N2109, N4673, N5509);
and AND4 (N6454, N6436, N4102, N5892, N4480);
and AND2 (N6455, N6447, N2398);
nor NOR4 (N6456, N6440, N2734, N5507, N726);
and AND4 (N6457, N6449, N4005, N4556, N2369);
nor NOR3 (N6458, N6452, N4843, N2479);
or OR2 (N6459, N6457, N2742);
not NOT1 (N6460, N6405);
and AND3 (N6461, N6456, N3565, N951);
and AND2 (N6462, N6430, N1924);
nand NAND3 (N6463, N6451, N51, N4278);
nand NAND2 (N6464, N6463, N5190);
nand NAND4 (N6465, N6458, N5131, N2428, N1892);
nand NAND2 (N6466, N6461, N5737);
and AND3 (N6467, N6464, N6070, N2861);
or OR2 (N6468, N6462, N4180);
nor NOR2 (N6469, N6455, N4983);
not NOT1 (N6470, N6460);
or OR3 (N6471, N6470, N2715, N2671);
buf BUF1 (N6472, N6468);
not NOT1 (N6473, N6453);
not NOT1 (N6474, N6454);
xor XOR2 (N6475, N6466, N2359);
and AND2 (N6476, N6422, N5009);
and AND2 (N6477, N6474, N5613);
nand NAND3 (N6478, N6465, N1289, N658);
buf BUF1 (N6479, N6477);
or OR4 (N6480, N6472, N415, N4277, N4839);
nand NAND3 (N6481, N6480, N2608, N96);
buf BUF1 (N6482, N6478);
not NOT1 (N6483, N6479);
buf BUF1 (N6484, N6471);
nor NOR3 (N6485, N6467, N2125, N3184);
or OR4 (N6486, N6459, N917, N6232, N4433);
nand NAND4 (N6487, N6469, N1287, N1726, N1229);
or OR2 (N6488, N6482, N4934);
and AND3 (N6489, N6484, N3719, N4310);
nand NAND3 (N6490, N6487, N3992, N4987);
nor NOR3 (N6491, N6475, N2937, N2418);
nand NAND4 (N6492, N6486, N6127, N5255, N4944);
or OR2 (N6493, N6490, N4024);
xor XOR2 (N6494, N6488, N368);
nor NOR2 (N6495, N6483, N3667);
or OR3 (N6496, N6491, N4722, N6482);
nand NAND3 (N6497, N6496, N4690, N5130);
buf BUF1 (N6498, N6489);
not NOT1 (N6499, N6476);
or OR4 (N6500, N6492, N3704, N3798, N414);
xor XOR2 (N6501, N6494, N1422);
or OR2 (N6502, N6497, N5368);
xor XOR2 (N6503, N6493, N5063);
xor XOR2 (N6504, N6498, N4871);
xor XOR2 (N6505, N6495, N2349);
or OR4 (N6506, N6500, N4932, N2257, N1536);
or OR2 (N6507, N6473, N6054);
or OR2 (N6508, N6504, N3641);
not NOT1 (N6509, N6501);
nor NOR2 (N6510, N6507, N1902);
and AND2 (N6511, N6481, N2314);
xor XOR2 (N6512, N6510, N5082);
and AND2 (N6513, N6512, N5121);
and AND3 (N6514, N6509, N2460, N4279);
buf BUF1 (N6515, N6499);
and AND2 (N6516, N6505, N2053);
nand NAND2 (N6517, N6511, N24);
not NOT1 (N6518, N6506);
and AND2 (N6519, N6503, N317);
nor NOR3 (N6520, N6515, N4402, N2422);
and AND4 (N6521, N6513, N3236, N4439, N3529);
buf BUF1 (N6522, N6517);
nor NOR2 (N6523, N6502, N6042);
and AND2 (N6524, N6485, N4685);
not NOT1 (N6525, N6508);
buf BUF1 (N6526, N6514);
nor NOR3 (N6527, N6518, N5998, N2658);
nand NAND4 (N6528, N6527, N1737, N1458, N4190);
or OR3 (N6529, N6528, N1614, N4140);
not NOT1 (N6530, N6526);
buf BUF1 (N6531, N6521);
not NOT1 (N6532, N6520);
or OR3 (N6533, N6523, N4408, N827);
and AND2 (N6534, N6516, N993);
or OR2 (N6535, N6530, N3233);
nand NAND3 (N6536, N6525, N160, N3663);
or OR2 (N6537, N6524, N5869);
or OR3 (N6538, N6535, N2563, N5577);
or OR4 (N6539, N6537, N5029, N1188, N5237);
and AND4 (N6540, N6531, N3295, N1857, N4499);
not NOT1 (N6541, N6532);
buf BUF1 (N6542, N6539);
not NOT1 (N6543, N6519);
xor XOR2 (N6544, N6540, N2991);
nor NOR4 (N6545, N6542, N3177, N5228, N4900);
not NOT1 (N6546, N6544);
nand NAND4 (N6547, N6533, N6392, N776, N5248);
not NOT1 (N6548, N6534);
and AND3 (N6549, N6545, N6471, N4748);
xor XOR2 (N6550, N6541, N2245);
nor NOR4 (N6551, N6546, N501, N658, N4341);
xor XOR2 (N6552, N6547, N2542);
not NOT1 (N6553, N6549);
nor NOR2 (N6554, N6543, N6121);
buf BUF1 (N6555, N6552);
buf BUF1 (N6556, N6536);
not NOT1 (N6557, N6554);
or OR4 (N6558, N6548, N3714, N2672, N2423);
xor XOR2 (N6559, N6556, N5815);
buf BUF1 (N6560, N6538);
xor XOR2 (N6561, N6553, N4440);
xor XOR2 (N6562, N6557, N5205);
buf BUF1 (N6563, N6522);
or OR2 (N6564, N6562, N4146);
not NOT1 (N6565, N6560);
nand NAND3 (N6566, N6561, N2199, N1140);
not NOT1 (N6567, N6550);
xor XOR2 (N6568, N6555, N2095);
nor NOR2 (N6569, N6564, N4610);
and AND2 (N6570, N6551, N4075);
xor XOR2 (N6571, N6559, N4531);
buf BUF1 (N6572, N6568);
buf BUF1 (N6573, N6563);
buf BUF1 (N6574, N6558);
or OR4 (N6575, N6565, N2601, N1413, N3766);
nand NAND2 (N6576, N6574, N6074);
buf BUF1 (N6577, N6571);
buf BUF1 (N6578, N6570);
not NOT1 (N6579, N6575);
xor XOR2 (N6580, N6573, N4983);
and AND3 (N6581, N6580, N1368, N324);
xor XOR2 (N6582, N6566, N5984);
or OR4 (N6583, N6578, N969, N4690, N1082);
not NOT1 (N6584, N6529);
xor XOR2 (N6585, N6579, N2490);
nand NAND3 (N6586, N6567, N2197, N3042);
or OR4 (N6587, N6572, N6252, N1877, N369);
nor NOR2 (N6588, N6576, N598);
not NOT1 (N6589, N6582);
buf BUF1 (N6590, N6577);
nor NOR4 (N6591, N6587, N4455, N4737, N4520);
and AND3 (N6592, N6584, N3214, N3587);
buf BUF1 (N6593, N6590);
buf BUF1 (N6594, N6589);
xor XOR2 (N6595, N6593, N5233);
not NOT1 (N6596, N6595);
nand NAND3 (N6597, N6592, N1633, N25);
buf BUF1 (N6598, N6569);
and AND4 (N6599, N6588, N6282, N4307, N1150);
buf BUF1 (N6600, N6598);
or OR3 (N6601, N6600, N3974, N1860);
not NOT1 (N6602, N6585);
xor XOR2 (N6603, N6586, N6144);
nor NOR4 (N6604, N6583, N682, N3129, N4178);
buf BUF1 (N6605, N6596);
and AND3 (N6606, N6599, N6420, N5087);
buf BUF1 (N6607, N6601);
nand NAND3 (N6608, N6606, N2058, N3024);
nor NOR2 (N6609, N6594, N3334);
nand NAND3 (N6610, N6591, N1139, N1267);
nor NOR4 (N6611, N6609, N636, N495, N5728);
or OR4 (N6612, N6581, N4117, N4719, N1714);
buf BUF1 (N6613, N6597);
nor NOR2 (N6614, N6612, N2753);
xor XOR2 (N6615, N6611, N3655);
and AND4 (N6616, N6610, N3570, N1484, N5541);
or OR4 (N6617, N6615, N2847, N2173, N3677);
nor NOR2 (N6618, N6617, N963);
xor XOR2 (N6619, N6613, N5574);
not NOT1 (N6620, N6619);
not NOT1 (N6621, N6618);
not NOT1 (N6622, N6602);
and AND3 (N6623, N6603, N1852, N916);
or OR4 (N6624, N6614, N4718, N1995, N4166);
and AND4 (N6625, N6621, N4125, N2390, N6155);
and AND3 (N6626, N6620, N6396, N4525);
not NOT1 (N6627, N6604);
not NOT1 (N6628, N6608);
nor NOR4 (N6629, N6628, N1632, N393, N3195);
and AND2 (N6630, N6627, N2671);
or OR4 (N6631, N6624, N4971, N948, N833);
or OR2 (N6632, N6607, N2173);
nand NAND2 (N6633, N6632, N797);
nor NOR3 (N6634, N6630, N1972, N3957);
or OR4 (N6635, N6616, N658, N5313, N6545);
and AND3 (N6636, N6623, N1152, N5972);
not NOT1 (N6637, N6634);
nand NAND4 (N6638, N6626, N4550, N4004, N5618);
nand NAND3 (N6639, N6636, N3900, N343);
buf BUF1 (N6640, N6631);
nand NAND2 (N6641, N6625, N1706);
not NOT1 (N6642, N6637);
xor XOR2 (N6643, N6639, N5397);
xor XOR2 (N6644, N6641, N6);
xor XOR2 (N6645, N6605, N5814);
xor XOR2 (N6646, N6640, N4458);
nor NOR2 (N6647, N6638, N5011);
not NOT1 (N6648, N6622);
xor XOR2 (N6649, N6644, N3489);
or OR4 (N6650, N6629, N5313, N3723, N2467);
nor NOR4 (N6651, N6650, N6136, N1186, N4183);
not NOT1 (N6652, N6649);
buf BUF1 (N6653, N6652);
nor NOR4 (N6654, N6642, N5137, N3757, N3757);
nand NAND2 (N6655, N6646, N595);
or OR3 (N6656, N6635, N4019, N4306);
nor NOR3 (N6657, N6647, N2938, N5469);
not NOT1 (N6658, N6656);
and AND4 (N6659, N6645, N3694, N6054, N1760);
nand NAND4 (N6660, N6658, N5041, N6529, N6442);
or OR4 (N6661, N6643, N2355, N2100, N1639);
not NOT1 (N6662, N6648);
and AND4 (N6663, N6654, N439, N5529, N3105);
not NOT1 (N6664, N6655);
nor NOR2 (N6665, N6633, N2518);
or OR2 (N6666, N6664, N639);
not NOT1 (N6667, N6660);
not NOT1 (N6668, N6662);
not NOT1 (N6669, N6665);
or OR2 (N6670, N6666, N5193);
xor XOR2 (N6671, N6669, N5639);
nand NAND4 (N6672, N6663, N368, N326, N5603);
or OR4 (N6673, N6659, N1141, N4517, N4038);
or OR2 (N6674, N6667, N4063);
not NOT1 (N6675, N6668);
nor NOR3 (N6676, N6661, N136, N777);
nand NAND3 (N6677, N6675, N4254, N3566);
not NOT1 (N6678, N6676);
buf BUF1 (N6679, N6678);
or OR2 (N6680, N6651, N6025);
nand NAND4 (N6681, N6671, N3132, N2358, N6375);
or OR4 (N6682, N6677, N1605, N3057, N6664);
nor NOR4 (N6683, N6680, N454, N463, N2286);
and AND3 (N6684, N6682, N4387, N1495);
buf BUF1 (N6685, N6673);
or OR3 (N6686, N6657, N4750, N4782);
not NOT1 (N6687, N6670);
or OR3 (N6688, N6674, N5182, N4842);
buf BUF1 (N6689, N6672);
and AND3 (N6690, N6653, N4540, N6131);
and AND4 (N6691, N6687, N2966, N1695, N69);
nor NOR4 (N6692, N6686, N3468, N3788, N6272);
nor NOR4 (N6693, N6692, N4079, N2132, N6136);
and AND2 (N6694, N6693, N71);
xor XOR2 (N6695, N6683, N2347);
or OR3 (N6696, N6684, N4996, N92);
and AND2 (N6697, N6688, N2751);
xor XOR2 (N6698, N6695, N4346);
nand NAND4 (N6699, N6697, N1990, N5502, N1796);
not NOT1 (N6700, N6690);
nand NAND2 (N6701, N6698, N1496);
not NOT1 (N6702, N6700);
xor XOR2 (N6703, N6694, N5111);
and AND4 (N6704, N6691, N1250, N5797, N4255);
buf BUF1 (N6705, N6679);
not NOT1 (N6706, N6703);
nand NAND4 (N6707, N6705, N3811, N4344, N5728);
not NOT1 (N6708, N6685);
nor NOR3 (N6709, N6699, N6095, N285);
buf BUF1 (N6710, N6681);
xor XOR2 (N6711, N6710, N1717);
buf BUF1 (N6712, N6704);
nor NOR2 (N6713, N6706, N852);
nor NOR4 (N6714, N6701, N5747, N2100, N3378);
xor XOR2 (N6715, N6696, N625);
nor NOR3 (N6716, N6714, N5688, N126);
xor XOR2 (N6717, N6708, N1375);
or OR2 (N6718, N6713, N5687);
or OR2 (N6719, N6711, N91);
or OR4 (N6720, N6715, N99, N5409, N5733);
not NOT1 (N6721, N6707);
xor XOR2 (N6722, N6716, N3254);
not NOT1 (N6723, N6709);
and AND3 (N6724, N6702, N2219, N6444);
or OR3 (N6725, N6689, N6111, N6572);
nor NOR3 (N6726, N6717, N2751, N6718);
xor XOR2 (N6727, N3033, N3631);
nand NAND3 (N6728, N6722, N4774, N6612);
xor XOR2 (N6729, N6720, N5045);
xor XOR2 (N6730, N6719, N4942);
not NOT1 (N6731, N6712);
or OR3 (N6732, N6725, N1439, N6357);
buf BUF1 (N6733, N6723);
nor NOR4 (N6734, N6726, N274, N965, N4086);
and AND2 (N6735, N6729, N779);
not NOT1 (N6736, N6721);
not NOT1 (N6737, N6728);
and AND2 (N6738, N6736, N5520);
and AND4 (N6739, N6738, N4148, N3319, N3399);
or OR3 (N6740, N6732, N4838, N5796);
and AND2 (N6741, N6737, N976);
nand NAND2 (N6742, N6724, N965);
or OR3 (N6743, N6740, N224, N6341);
nand NAND4 (N6744, N6735, N2003, N2714, N6662);
and AND2 (N6745, N6727, N4066);
xor XOR2 (N6746, N6730, N1661);
nand NAND2 (N6747, N6733, N4637);
xor XOR2 (N6748, N6745, N3896);
nor NOR4 (N6749, N6742, N1627, N3020, N1216);
nand NAND4 (N6750, N6744, N6301, N1757, N1004);
not NOT1 (N6751, N6750);
not NOT1 (N6752, N6747);
not NOT1 (N6753, N6741);
or OR4 (N6754, N6752, N983, N80, N5093);
xor XOR2 (N6755, N6739, N3689);
nor NOR4 (N6756, N6755, N388, N679, N4996);
not NOT1 (N6757, N6754);
nand NAND3 (N6758, N6753, N1008, N3336);
not NOT1 (N6759, N6756);
xor XOR2 (N6760, N6748, N1645);
nand NAND2 (N6761, N6731, N2680);
nor NOR3 (N6762, N6761, N3156, N1518);
not NOT1 (N6763, N6760);
buf BUF1 (N6764, N6746);
and AND3 (N6765, N6763, N4528, N5894);
and AND3 (N6766, N6734, N1053, N3935);
nor NOR2 (N6767, N6751, N1263);
and AND2 (N6768, N6765, N730);
not NOT1 (N6769, N6749);
or OR3 (N6770, N6767, N790, N6478);
or OR3 (N6771, N6764, N2573, N6240);
xor XOR2 (N6772, N6768, N2448);
buf BUF1 (N6773, N6743);
nor NOR2 (N6774, N6759, N5816);
or OR3 (N6775, N6773, N4870, N3435);
buf BUF1 (N6776, N6774);
not NOT1 (N6777, N6775);
not NOT1 (N6778, N6777);
nand NAND4 (N6779, N6776, N3973, N794, N1215);
not NOT1 (N6780, N6770);
nand NAND4 (N6781, N6772, N2683, N439, N1277);
or OR3 (N6782, N6778, N2160, N1578);
buf BUF1 (N6783, N6782);
or OR2 (N6784, N6783, N3661);
nor NOR2 (N6785, N6784, N2607);
nor NOR4 (N6786, N6779, N3886, N1260, N4622);
nand NAND2 (N6787, N6762, N5961);
nor NOR2 (N6788, N6781, N5933);
not NOT1 (N6789, N6780);
or OR3 (N6790, N6786, N2178, N4783);
nor NOR4 (N6791, N6790, N6368, N2388, N5081);
not NOT1 (N6792, N6758);
nand NAND2 (N6793, N6787, N1820);
not NOT1 (N6794, N6788);
xor XOR2 (N6795, N6791, N5259);
nand NAND3 (N6796, N6757, N1622, N133);
buf BUF1 (N6797, N6793);
xor XOR2 (N6798, N6795, N3638);
nand NAND4 (N6799, N6794, N5572, N820, N354);
or OR2 (N6800, N6766, N6421);
nand NAND3 (N6801, N6796, N6759, N1075);
not NOT1 (N6802, N6800);
nand NAND4 (N6803, N6797, N649, N3336, N433);
xor XOR2 (N6804, N6798, N5699);
not NOT1 (N6805, N6769);
or OR3 (N6806, N6801, N2059, N315);
not NOT1 (N6807, N6804);
and AND4 (N6808, N6806, N1887, N4859, N1184);
nor NOR4 (N6809, N6789, N6148, N783, N2120);
buf BUF1 (N6810, N6809);
buf BUF1 (N6811, N6771);
nor NOR4 (N6812, N6785, N2361, N4927, N1222);
xor XOR2 (N6813, N6802, N6396);
or OR4 (N6814, N6799, N5514, N3657, N4556);
nand NAND4 (N6815, N6808, N6070, N268, N2180);
not NOT1 (N6816, N6810);
not NOT1 (N6817, N6814);
xor XOR2 (N6818, N6807, N5537);
or OR3 (N6819, N6792, N3406, N398);
or OR4 (N6820, N6805, N1201, N1014, N2749);
not NOT1 (N6821, N6816);
nor NOR2 (N6822, N6821, N1540);
nand NAND2 (N6823, N6812, N3065);
or OR3 (N6824, N6813, N5895, N2831);
buf BUF1 (N6825, N6815);
xor XOR2 (N6826, N6819, N4898);
buf BUF1 (N6827, N6822);
nor NOR4 (N6828, N6824, N5263, N1948, N3968);
nor NOR4 (N6829, N6825, N3111, N5488, N2053);
and AND3 (N6830, N6817, N3039, N5905);
xor XOR2 (N6831, N6830, N3215);
not NOT1 (N6832, N6811);
nand NAND2 (N6833, N6818, N2248);
not NOT1 (N6834, N6828);
or OR3 (N6835, N6827, N2902, N6792);
xor XOR2 (N6836, N6829, N5332);
and AND2 (N6837, N6834, N2975);
or OR2 (N6838, N6836, N850);
xor XOR2 (N6839, N6826, N3785);
not NOT1 (N6840, N6832);
not NOT1 (N6841, N6839);
and AND4 (N6842, N6840, N5966, N2892, N4285);
nand NAND3 (N6843, N6835, N5425, N496);
not NOT1 (N6844, N6823);
buf BUF1 (N6845, N6838);
or OR4 (N6846, N6833, N3626, N6343, N6755);
buf BUF1 (N6847, N6837);
buf BUF1 (N6848, N6842);
xor XOR2 (N6849, N6831, N6498);
nand NAND3 (N6850, N6847, N6297, N5716);
buf BUF1 (N6851, N6803);
nand NAND3 (N6852, N6851, N373, N2795);
xor XOR2 (N6853, N6820, N2642);
xor XOR2 (N6854, N6845, N1712);
nand NAND4 (N6855, N6853, N2579, N4632, N5971);
or OR2 (N6856, N6846, N107);
nor NOR4 (N6857, N6855, N3147, N3936, N3537);
nand NAND3 (N6858, N6852, N3105, N6615);
nor NOR3 (N6859, N6857, N6240, N2109);
nand NAND3 (N6860, N6849, N5905, N1947);
nor NOR2 (N6861, N6850, N6410);
or OR2 (N6862, N6856, N5919);
and AND4 (N6863, N6843, N1280, N5410, N2695);
or OR3 (N6864, N6863, N5627, N5118);
buf BUF1 (N6865, N6862);
or OR3 (N6866, N6860, N3931, N5338);
buf BUF1 (N6867, N6858);
and AND3 (N6868, N6865, N943, N1491);
nor NOR3 (N6869, N6859, N3648, N3513);
buf BUF1 (N6870, N6841);
nor NOR2 (N6871, N6848, N4178);
nor NOR3 (N6872, N6870, N1821, N1014);
nor NOR3 (N6873, N6871, N2670, N3952);
nand NAND2 (N6874, N6864, N1021);
not NOT1 (N6875, N6844);
nor NOR2 (N6876, N6866, N6112);
buf BUF1 (N6877, N6867);
and AND2 (N6878, N6854, N1092);
or OR3 (N6879, N6868, N1165, N5083);
nor NOR3 (N6880, N6877, N523, N1254);
buf BUF1 (N6881, N6875);
nand NAND4 (N6882, N6878, N6649, N5899, N2867);
nand NAND2 (N6883, N6869, N2745);
nand NAND3 (N6884, N6882, N4786, N5026);
nor NOR2 (N6885, N6883, N337);
xor XOR2 (N6886, N6884, N6122);
nor NOR4 (N6887, N6876, N4762, N3490, N5061);
nor NOR2 (N6888, N6879, N6544);
or OR2 (N6889, N6861, N2881);
and AND3 (N6890, N6887, N2988, N3359);
xor XOR2 (N6891, N6880, N2671);
xor XOR2 (N6892, N6885, N4369);
nand NAND2 (N6893, N6890, N6001);
nand NAND4 (N6894, N6873, N2163, N223, N3623);
nor NOR2 (N6895, N6888, N3369);
xor XOR2 (N6896, N6892, N2554);
xor XOR2 (N6897, N6886, N5475);
and AND3 (N6898, N6891, N3729, N1344);
nand NAND2 (N6899, N6898, N3997);
buf BUF1 (N6900, N6881);
buf BUF1 (N6901, N6897);
nand NAND2 (N6902, N6894, N3223);
or OR2 (N6903, N6893, N5878);
nand NAND4 (N6904, N6902, N2788, N5645, N767);
or OR3 (N6905, N6904, N6006, N1913);
nand NAND3 (N6906, N6901, N1634, N3510);
nor NOR4 (N6907, N6906, N3389, N5646, N5121);
nor NOR3 (N6908, N6895, N5916, N4678);
nor NOR3 (N6909, N6872, N6321, N766);
nor NOR4 (N6910, N6908, N2528, N2165, N810);
not NOT1 (N6911, N6910);
or OR3 (N6912, N6874, N3385, N4467);
or OR4 (N6913, N6912, N45, N1597, N3231);
not NOT1 (N6914, N6889);
or OR2 (N6915, N6914, N6699);
or OR4 (N6916, N6915, N250, N6094, N1594);
and AND4 (N6917, N6899, N1273, N2572, N5376);
nand NAND2 (N6918, N6896, N6389);
xor XOR2 (N6919, N6900, N1252);
nor NOR4 (N6920, N6913, N2175, N6731, N5971);
buf BUF1 (N6921, N6907);
nand NAND3 (N6922, N6905, N6055, N6119);
nand NAND2 (N6923, N6919, N3360);
nand NAND2 (N6924, N6922, N2840);
xor XOR2 (N6925, N6917, N658);
xor XOR2 (N6926, N6924, N2978);
nor NOR4 (N6927, N6926, N6173, N354, N3598);
xor XOR2 (N6928, N6920, N1049);
or OR4 (N6929, N6918, N6160, N4892, N274);
buf BUF1 (N6930, N6927);
nand NAND4 (N6931, N6923, N4786, N937, N2057);
or OR4 (N6932, N6921, N854, N3676, N4635);
not NOT1 (N6933, N6911);
and AND3 (N6934, N6909, N4945, N1897);
not NOT1 (N6935, N6930);
buf BUF1 (N6936, N6933);
and AND4 (N6937, N6928, N3600, N2753, N6671);
nand NAND4 (N6938, N6936, N512, N2333, N2376);
nand NAND3 (N6939, N6935, N6240, N2341);
nand NAND3 (N6940, N6903, N3161, N3785);
nand NAND2 (N6941, N6929, N4642);
not NOT1 (N6942, N6941);
and AND2 (N6943, N6938, N5362);
not NOT1 (N6944, N6932);
and AND3 (N6945, N6916, N501, N425);
xor XOR2 (N6946, N6945, N3257);
and AND4 (N6947, N6943, N6460, N1964, N2165);
nand NAND3 (N6948, N6925, N6236, N2199);
nand NAND2 (N6949, N6942, N2599);
and AND3 (N6950, N6944, N3510, N1536);
or OR3 (N6951, N6940, N5498, N350);
or OR3 (N6952, N6949, N2366, N5311);
xor XOR2 (N6953, N6931, N126);
nor NOR4 (N6954, N6951, N920, N6581, N3487);
nor NOR2 (N6955, N6952, N6228);
xor XOR2 (N6956, N6946, N2091);
buf BUF1 (N6957, N6953);
nor NOR2 (N6958, N6934, N4003);
not NOT1 (N6959, N6955);
not NOT1 (N6960, N6948);
nor NOR4 (N6961, N6947, N1422, N3730, N45);
and AND4 (N6962, N6956, N6154, N383, N3466);
nor NOR4 (N6963, N6959, N6316, N772, N2838);
not NOT1 (N6964, N6963);
nand NAND3 (N6965, N6950, N4558, N2743);
or OR2 (N6966, N6957, N3326);
not NOT1 (N6967, N6937);
and AND4 (N6968, N6958, N2361, N5071, N3208);
or OR4 (N6969, N6964, N2909, N210, N6237);
buf BUF1 (N6970, N6967);
xor XOR2 (N6971, N6960, N6188);
or OR2 (N6972, N6966, N5115);
xor XOR2 (N6973, N6965, N2309);
nor NOR4 (N6974, N6971, N5030, N3140, N137);
not NOT1 (N6975, N6968);
xor XOR2 (N6976, N6973, N2165);
nor NOR4 (N6977, N6954, N4733, N994, N5041);
nor NOR2 (N6978, N6974, N2027);
or OR4 (N6979, N6978, N1722, N3361, N358);
nand NAND2 (N6980, N6975, N4589);
buf BUF1 (N6981, N6977);
or OR4 (N6982, N6979, N694, N1710, N6037);
and AND2 (N6983, N6980, N4476);
nand NAND2 (N6984, N6981, N2039);
or OR3 (N6985, N6984, N89, N548);
nand NAND3 (N6986, N6976, N284, N2732);
not NOT1 (N6987, N6982);
not NOT1 (N6988, N6962);
nand NAND2 (N6989, N6969, N5151);
buf BUF1 (N6990, N6986);
buf BUF1 (N6991, N6985);
nor NOR3 (N6992, N6987, N3020, N2876);
nor NOR3 (N6993, N6983, N6137, N1927);
buf BUF1 (N6994, N6991);
buf BUF1 (N6995, N6961);
or OR2 (N6996, N6994, N6668);
and AND4 (N6997, N6996, N2377, N1990, N4494);
nand NAND3 (N6998, N6995, N6758, N3145);
buf BUF1 (N6999, N6997);
nor NOR3 (N7000, N6970, N3639, N4105);
nor NOR3 (N7001, N6989, N1945, N2523);
nor NOR2 (N7002, N6992, N3714);
xor XOR2 (N7003, N6972, N1483);
nand NAND3 (N7004, N7002, N4547, N483);
buf BUF1 (N7005, N6988);
nor NOR3 (N7006, N7004, N2102, N1309);
nand NAND2 (N7007, N6993, N486);
nor NOR4 (N7008, N6939, N6937, N5560, N4734);
xor XOR2 (N7009, N7008, N4903);
nor NOR2 (N7010, N7003, N6066);
or OR3 (N7011, N7000, N3376, N877);
nand NAND2 (N7012, N7009, N715);
nand NAND2 (N7013, N7012, N1680);
and AND2 (N7014, N6998, N6035);
buf BUF1 (N7015, N7007);
or OR2 (N7016, N7005, N2262);
not NOT1 (N7017, N6999);
or OR4 (N7018, N6990, N6423, N3471, N1548);
or OR2 (N7019, N7017, N3892);
nor NOR3 (N7020, N7001, N6432, N6712);
not NOT1 (N7021, N7014);
or OR4 (N7022, N7018, N958, N3617, N2287);
nand NAND3 (N7023, N7011, N4969, N973);
and AND3 (N7024, N7016, N245, N2428);
or OR4 (N7025, N7006, N6743, N1146, N2113);
xor XOR2 (N7026, N7021, N1324);
xor XOR2 (N7027, N7020, N3950);
or OR3 (N7028, N7015, N6374, N1991);
buf BUF1 (N7029, N7019);
not NOT1 (N7030, N7026);
and AND2 (N7031, N7028, N6310);
not NOT1 (N7032, N7030);
xor XOR2 (N7033, N7027, N35);
or OR3 (N7034, N7033, N5872, N3531);
and AND4 (N7035, N7010, N5863, N3457, N5652);
or OR2 (N7036, N7013, N2486);
buf BUF1 (N7037, N7036);
or OR3 (N7038, N7034, N4310, N6152);
nand NAND4 (N7039, N7038, N886, N2055, N6749);
not NOT1 (N7040, N7025);
buf BUF1 (N7041, N7035);
not NOT1 (N7042, N7037);
xor XOR2 (N7043, N7040, N1574);
nand NAND3 (N7044, N7039, N1446, N1844);
not NOT1 (N7045, N7041);
nor NOR3 (N7046, N7029, N3607, N1319);
nor NOR3 (N7047, N7045, N6102, N3437);
or OR2 (N7048, N7024, N3981);
and AND4 (N7049, N7023, N1461, N6782, N6090);
not NOT1 (N7050, N7049);
or OR4 (N7051, N7043, N5742, N3871, N1629);
buf BUF1 (N7052, N7050);
buf BUF1 (N7053, N7032);
buf BUF1 (N7054, N7048);
not NOT1 (N7055, N7046);
not NOT1 (N7056, N7044);
nand NAND3 (N7057, N7052, N6785, N2092);
and AND4 (N7058, N7055, N2419, N3944, N229);
nor NOR4 (N7059, N7047, N4616, N4408, N4467);
or OR2 (N7060, N7022, N3939);
nor NOR2 (N7061, N7058, N941);
buf BUF1 (N7062, N7059);
or OR4 (N7063, N7060, N3673, N4941, N684);
and AND3 (N7064, N7063, N4050, N2214);
and AND2 (N7065, N7031, N3202);
or OR4 (N7066, N7065, N3071, N6330, N5752);
and AND2 (N7067, N7062, N904);
nor NOR3 (N7068, N7064, N3142, N4885);
and AND4 (N7069, N7067, N4883, N2854, N158);
xor XOR2 (N7070, N7057, N3203);
not NOT1 (N7071, N7042);
or OR4 (N7072, N7054, N5206, N778, N5315);
xor XOR2 (N7073, N7068, N108);
buf BUF1 (N7074, N7066);
not NOT1 (N7075, N7073);
nand NAND3 (N7076, N7070, N1599, N6291);
nor NOR3 (N7077, N7075, N717, N6030);
buf BUF1 (N7078, N7076);
or OR3 (N7079, N7078, N2909, N1267);
buf BUF1 (N7080, N7056);
not NOT1 (N7081, N7079);
nand NAND3 (N7082, N7072, N6267, N1752);
buf BUF1 (N7083, N7082);
not NOT1 (N7084, N7069);
nor NOR4 (N7085, N7080, N2368, N2242, N4257);
or OR4 (N7086, N7084, N4106, N6072, N565);
buf BUF1 (N7087, N7051);
and AND4 (N7088, N7087, N3769, N1970, N4626);
buf BUF1 (N7089, N7061);
buf BUF1 (N7090, N7071);
nand NAND3 (N7091, N7088, N3971, N3133);
nand NAND4 (N7092, N7081, N4228, N4229, N5);
or OR2 (N7093, N7089, N1093);
xor XOR2 (N7094, N7093, N5724);
or OR2 (N7095, N7092, N1968);
nand NAND4 (N7096, N7083, N146, N2254, N3572);
buf BUF1 (N7097, N7091);
and AND3 (N7098, N7086, N388, N715);
xor XOR2 (N7099, N7098, N6347);
not NOT1 (N7100, N7090);
or OR3 (N7101, N7096, N2001, N585);
or OR3 (N7102, N7053, N883, N4852);
buf BUF1 (N7103, N7100);
not NOT1 (N7104, N7085);
xor XOR2 (N7105, N7103, N6057);
and AND2 (N7106, N7101, N3141);
xor XOR2 (N7107, N7102, N5912);
buf BUF1 (N7108, N7074);
and AND3 (N7109, N7099, N6655, N6024);
or OR3 (N7110, N7095, N3607, N2855);
and AND2 (N7111, N7094, N5090);
not NOT1 (N7112, N7111);
xor XOR2 (N7113, N7112, N4561);
buf BUF1 (N7114, N7110);
buf BUF1 (N7115, N7097);
xor XOR2 (N7116, N7113, N2067);
buf BUF1 (N7117, N7105);
xor XOR2 (N7118, N7114, N5540);
nor NOR2 (N7119, N7118, N1744);
nand NAND2 (N7120, N7107, N579);
nor NOR4 (N7121, N7115, N2835, N2368, N3665);
and AND2 (N7122, N7108, N6621);
not NOT1 (N7123, N7077);
not NOT1 (N7124, N7104);
buf BUF1 (N7125, N7106);
not NOT1 (N7126, N7123);
xor XOR2 (N7127, N7109, N6371);
not NOT1 (N7128, N7120);
buf BUF1 (N7129, N7116);
nand NAND3 (N7130, N7122, N2939, N6426);
buf BUF1 (N7131, N7129);
or OR2 (N7132, N7128, N3284);
and AND2 (N7133, N7126, N6292);
not NOT1 (N7134, N7124);
nor NOR3 (N7135, N7127, N1171, N881);
and AND4 (N7136, N7135, N1183, N4610, N4144);
nor NOR2 (N7137, N7136, N6215);
xor XOR2 (N7138, N7132, N5472);
nor NOR2 (N7139, N7137, N6148);
nor NOR2 (N7140, N7131, N2177);
nand NAND4 (N7141, N7138, N2043, N1255, N6986);
or OR3 (N7142, N7141, N341, N5317);
xor XOR2 (N7143, N7130, N6009);
xor XOR2 (N7144, N7119, N1447);
and AND2 (N7145, N7117, N4299);
and AND4 (N7146, N7134, N6692, N125, N3455);
xor XOR2 (N7147, N7144, N1586);
xor XOR2 (N7148, N7133, N3018);
not NOT1 (N7149, N7125);
and AND4 (N7150, N7139, N4039, N3575, N4393);
or OR3 (N7151, N7143, N4719, N2143);
not NOT1 (N7152, N7145);
nand NAND2 (N7153, N7142, N451);
and AND4 (N7154, N7146, N5460, N5381, N4570);
not NOT1 (N7155, N7149);
nand NAND2 (N7156, N7153, N4276);
not NOT1 (N7157, N7121);
nand NAND3 (N7158, N7140, N1988, N3062);
nor NOR3 (N7159, N7150, N3734, N3165);
and AND3 (N7160, N7157, N4651, N7117);
nor NOR3 (N7161, N7152, N3995, N1677);
buf BUF1 (N7162, N7160);
nand NAND3 (N7163, N7154, N6025, N6867);
and AND4 (N7164, N7158, N817, N1215, N1098);
nand NAND2 (N7165, N7151, N4471);
not NOT1 (N7166, N7155);
buf BUF1 (N7167, N7161);
xor XOR2 (N7168, N7165, N3689);
or OR2 (N7169, N7163, N5202);
nand NAND4 (N7170, N7166, N1096, N5156, N2988);
buf BUF1 (N7171, N7162);
nand NAND4 (N7172, N7169, N2851, N2435, N1317);
xor XOR2 (N7173, N7147, N6172);
or OR2 (N7174, N7156, N2437);
buf BUF1 (N7175, N7168);
and AND2 (N7176, N7174, N4637);
buf BUF1 (N7177, N7172);
nor NOR3 (N7178, N7176, N574, N3089);
xor XOR2 (N7179, N7164, N5044);
nor NOR2 (N7180, N7178, N3151);
nand NAND3 (N7181, N7170, N1995, N966);
buf BUF1 (N7182, N7177);
not NOT1 (N7183, N7167);
and AND2 (N7184, N7181, N5429);
buf BUF1 (N7185, N7148);
nor NOR2 (N7186, N7173, N3555);
not NOT1 (N7187, N7186);
not NOT1 (N7188, N7171);
nor NOR3 (N7189, N7180, N6713, N5512);
and AND3 (N7190, N7187, N2904, N3913);
xor XOR2 (N7191, N7184, N7148);
nor NOR4 (N7192, N7179, N5090, N6362, N3530);
or OR2 (N7193, N7183, N1183);
nand NAND3 (N7194, N7189, N3239, N3865);
or OR3 (N7195, N7194, N3907, N775);
not NOT1 (N7196, N7185);
xor XOR2 (N7197, N7192, N2598);
buf BUF1 (N7198, N7182);
not NOT1 (N7199, N7196);
and AND2 (N7200, N7197, N4679);
nor NOR3 (N7201, N7198, N3981, N6650);
and AND2 (N7202, N7193, N3084);
xor XOR2 (N7203, N7191, N6184);
not NOT1 (N7204, N7159);
or OR4 (N7205, N7199, N2326, N6371, N5223);
buf BUF1 (N7206, N7190);
xor XOR2 (N7207, N7204, N5282);
buf BUF1 (N7208, N7195);
or OR4 (N7209, N7207, N5739, N4066, N2036);
xor XOR2 (N7210, N7205, N3245);
not NOT1 (N7211, N7188);
buf BUF1 (N7212, N7200);
xor XOR2 (N7213, N7203, N4786);
not NOT1 (N7214, N7175);
not NOT1 (N7215, N7209);
not NOT1 (N7216, N7212);
nand NAND3 (N7217, N7211, N3502, N4220);
buf BUF1 (N7218, N7201);
not NOT1 (N7219, N7213);
not NOT1 (N7220, N7208);
nand NAND4 (N7221, N7220, N3065, N5610, N5875);
xor XOR2 (N7222, N7221, N3518);
and AND2 (N7223, N7218, N7096);
nor NOR3 (N7224, N7219, N7089, N2659);
xor XOR2 (N7225, N7215, N1672);
buf BUF1 (N7226, N7216);
xor XOR2 (N7227, N7210, N4574);
not NOT1 (N7228, N7222);
xor XOR2 (N7229, N7202, N1892);
nor NOR4 (N7230, N7226, N1006, N243, N4350);
nand NAND3 (N7231, N7228, N2428, N3559);
buf BUF1 (N7232, N7229);
nand NAND3 (N7233, N7230, N419, N5445);
or OR4 (N7234, N7227, N5044, N4012, N3980);
nand NAND3 (N7235, N7214, N5157, N1262);
xor XOR2 (N7236, N7235, N6182);
not NOT1 (N7237, N7206);
or OR2 (N7238, N7224, N1259);
or OR2 (N7239, N7234, N2034);
or OR3 (N7240, N7217, N7225, N6202);
nand NAND3 (N7241, N5172, N5447, N5452);
nor NOR2 (N7242, N7231, N4637);
xor XOR2 (N7243, N7238, N3670);
xor XOR2 (N7244, N7243, N4967);
and AND4 (N7245, N7237, N782, N5865, N641);
and AND2 (N7246, N7242, N1396);
not NOT1 (N7247, N7246);
and AND2 (N7248, N7233, N1821);
buf BUF1 (N7249, N7236);
not NOT1 (N7250, N7232);
buf BUF1 (N7251, N7247);
nor NOR2 (N7252, N7248, N4528);
nor NOR3 (N7253, N7241, N5322, N1553);
buf BUF1 (N7254, N7245);
xor XOR2 (N7255, N7251, N5096);
and AND3 (N7256, N7252, N5806, N252);
not NOT1 (N7257, N7244);
nand NAND3 (N7258, N7254, N5861, N3564);
not NOT1 (N7259, N7239);
not NOT1 (N7260, N7253);
nand NAND4 (N7261, N7249, N5948, N3159, N6556);
or OR3 (N7262, N7255, N255, N4030);
or OR3 (N7263, N7262, N2752, N5739);
not NOT1 (N7264, N7260);
nand NAND2 (N7265, N7258, N3230);
xor XOR2 (N7266, N7263, N670);
and AND2 (N7267, N7250, N4212);
nand NAND2 (N7268, N7267, N1806);
nor NOR2 (N7269, N7256, N4843);
xor XOR2 (N7270, N7268, N1872);
buf BUF1 (N7271, N7257);
buf BUF1 (N7272, N7261);
or OR2 (N7273, N7265, N3760);
not NOT1 (N7274, N7264);
buf BUF1 (N7275, N7273);
buf BUF1 (N7276, N7275);
buf BUF1 (N7277, N7274);
and AND3 (N7278, N7276, N3297, N3038);
xor XOR2 (N7279, N7272, N6911);
not NOT1 (N7280, N7271);
nand NAND3 (N7281, N7269, N5028, N965);
or OR4 (N7282, N7223, N3002, N454, N2680);
and AND3 (N7283, N7282, N2293, N544);
xor XOR2 (N7284, N7259, N1276);
xor XOR2 (N7285, N7277, N5452);
nor NOR3 (N7286, N7266, N4391, N1959);
nor NOR2 (N7287, N7283, N4378);
buf BUF1 (N7288, N7281);
xor XOR2 (N7289, N7240, N3399);
xor XOR2 (N7290, N7287, N2166);
buf BUF1 (N7291, N7286);
nand NAND4 (N7292, N7285, N5388, N918, N4374);
and AND3 (N7293, N7292, N3340, N5326);
buf BUF1 (N7294, N7278);
nor NOR2 (N7295, N7293, N2027);
buf BUF1 (N7296, N7289);
xor XOR2 (N7297, N7290, N5691);
nor NOR3 (N7298, N7294, N5986, N4187);
and AND4 (N7299, N7296, N6710, N1294, N4562);
and AND2 (N7300, N7291, N3332);
xor XOR2 (N7301, N7297, N4469);
buf BUF1 (N7302, N7279);
xor XOR2 (N7303, N7298, N4398);
nand NAND2 (N7304, N7299, N5900);
and AND4 (N7305, N7303, N2235, N111, N5383);
nor NOR4 (N7306, N7300, N7195, N6235, N5880);
and AND2 (N7307, N7306, N305);
or OR2 (N7308, N7280, N4187);
nand NAND3 (N7309, N7295, N6265, N2598);
xor XOR2 (N7310, N7307, N2617);
or OR3 (N7311, N7302, N7176, N2390);
buf BUF1 (N7312, N7310);
xor XOR2 (N7313, N7304, N1054);
xor XOR2 (N7314, N7301, N5214);
nor NOR4 (N7315, N7309, N1910, N1662, N4963);
and AND4 (N7316, N7284, N1429, N4444, N7086);
not NOT1 (N7317, N7270);
nor NOR3 (N7318, N7308, N572, N7284);
or OR3 (N7319, N7305, N4208, N5522);
xor XOR2 (N7320, N7313, N341);
nor NOR4 (N7321, N7288, N7003, N6779, N466);
and AND2 (N7322, N7320, N4399);
nor NOR3 (N7323, N7315, N883, N6028);
xor XOR2 (N7324, N7312, N6737);
nand NAND3 (N7325, N7316, N4815, N1176);
xor XOR2 (N7326, N7322, N6879);
buf BUF1 (N7327, N7324);
nand NAND2 (N7328, N7319, N6529);
buf BUF1 (N7329, N7323);
buf BUF1 (N7330, N7328);
not NOT1 (N7331, N7325);
nor NOR4 (N7332, N7326, N106, N4127, N1004);
or OR4 (N7333, N7318, N573, N4891, N2221);
buf BUF1 (N7334, N7314);
or OR4 (N7335, N7327, N6134, N302, N3203);
nand NAND4 (N7336, N7331, N6756, N713, N2703);
and AND4 (N7337, N7332, N1237, N3465, N7098);
buf BUF1 (N7338, N7333);
or OR3 (N7339, N7334, N5954, N3958);
not NOT1 (N7340, N7317);
xor XOR2 (N7341, N7336, N4778);
buf BUF1 (N7342, N7335);
or OR3 (N7343, N7311, N6049, N2191);
or OR3 (N7344, N7341, N2096, N777);
or OR2 (N7345, N7340, N3530);
nand NAND2 (N7346, N7343, N5868);
or OR4 (N7347, N7346, N2275, N6696, N2961);
buf BUF1 (N7348, N7338);
not NOT1 (N7349, N7348);
buf BUF1 (N7350, N7344);
or OR2 (N7351, N7345, N5947);
nand NAND2 (N7352, N7339, N6205);
nand NAND2 (N7353, N7337, N1157);
and AND4 (N7354, N7321, N2622, N96, N6070);
xor XOR2 (N7355, N7347, N4422);
nand NAND2 (N7356, N7353, N1324);
nor NOR3 (N7357, N7355, N956, N4292);
and AND2 (N7358, N7349, N2113);
or OR4 (N7359, N7350, N603, N2592, N413);
and AND2 (N7360, N7354, N2044);
xor XOR2 (N7361, N7358, N257);
and AND4 (N7362, N7359, N155, N5472, N2715);
buf BUF1 (N7363, N7352);
buf BUF1 (N7364, N7356);
nor NOR3 (N7365, N7330, N6, N5651);
or OR3 (N7366, N7364, N347, N6024);
nand NAND2 (N7367, N7342, N6130);
and AND2 (N7368, N7367, N6698);
xor XOR2 (N7369, N7360, N2795);
nand NAND3 (N7370, N7351, N6945, N2822);
buf BUF1 (N7371, N7363);
not NOT1 (N7372, N7368);
nor NOR2 (N7373, N7366, N855);
and AND2 (N7374, N7370, N2051);
or OR4 (N7375, N7329, N4175, N2573, N5146);
not NOT1 (N7376, N7371);
xor XOR2 (N7377, N7361, N4708);
or OR3 (N7378, N7365, N6182, N3734);
nand NAND4 (N7379, N7377, N6593, N732, N7223);
xor XOR2 (N7380, N7372, N7209);
or OR3 (N7381, N7369, N3649, N5686);
nor NOR2 (N7382, N7380, N4588);
buf BUF1 (N7383, N7357);
not NOT1 (N7384, N7381);
nor NOR3 (N7385, N7379, N2800, N2093);
nand NAND2 (N7386, N7378, N3972);
or OR2 (N7387, N7373, N7380);
and AND3 (N7388, N7384, N4531, N1590);
or OR4 (N7389, N7385, N6667, N3519, N2224);
buf BUF1 (N7390, N7387);
nand NAND4 (N7391, N7388, N1223, N5710, N2240);
buf BUF1 (N7392, N7389);
nor NOR2 (N7393, N7391, N5044);
xor XOR2 (N7394, N7374, N915);
xor XOR2 (N7395, N7362, N2600);
or OR4 (N7396, N7395, N2921, N7295, N2380);
buf BUF1 (N7397, N7376);
not NOT1 (N7398, N7390);
nand NAND4 (N7399, N7396, N1226, N674, N4118);
or OR3 (N7400, N7375, N5322, N1173);
buf BUF1 (N7401, N7386);
buf BUF1 (N7402, N7392);
or OR4 (N7403, N7400, N5319, N4942, N1618);
xor XOR2 (N7404, N7397, N2130);
not NOT1 (N7405, N7403);
and AND3 (N7406, N7402, N4496, N6720);
nand NAND2 (N7407, N7404, N711);
nor NOR3 (N7408, N7406, N1202, N2926);
xor XOR2 (N7409, N7382, N3256);
nand NAND2 (N7410, N7409, N5124);
not NOT1 (N7411, N7407);
xor XOR2 (N7412, N7399, N5486);
nor NOR2 (N7413, N7394, N6390);
buf BUF1 (N7414, N7412);
nor NOR3 (N7415, N7413, N3864, N5148);
and AND3 (N7416, N7410, N763, N2995);
and AND3 (N7417, N7414, N7083, N3915);
xor XOR2 (N7418, N7415, N2581);
xor XOR2 (N7419, N7418, N3506);
buf BUF1 (N7420, N7411);
nand NAND4 (N7421, N7420, N2471, N6275, N4689);
xor XOR2 (N7422, N7383, N4302);
buf BUF1 (N7423, N7398);
buf BUF1 (N7424, N7423);
or OR2 (N7425, N7421, N880);
buf BUF1 (N7426, N7417);
buf BUF1 (N7427, N7422);
and AND2 (N7428, N7401, N4393);
nor NOR3 (N7429, N7419, N4237, N6775);
or OR2 (N7430, N7426, N5927);
or OR4 (N7431, N7393, N3744, N7070, N5379);
nor NOR3 (N7432, N7430, N5240, N2878);
not NOT1 (N7433, N7427);
or OR2 (N7434, N7431, N3689);
or OR3 (N7435, N7408, N2942, N3454);
buf BUF1 (N7436, N7428);
xor XOR2 (N7437, N7433, N3912);
nor NOR3 (N7438, N7437, N2550, N1549);
not NOT1 (N7439, N7416);
xor XOR2 (N7440, N7439, N2635);
not NOT1 (N7441, N7435);
not NOT1 (N7442, N7438);
xor XOR2 (N7443, N7441, N4071);
or OR2 (N7444, N7436, N1494);
xor XOR2 (N7445, N7443, N5833);
nand NAND4 (N7446, N7442, N4030, N2155, N5421);
and AND2 (N7447, N7444, N1943);
buf BUF1 (N7448, N7405);
or OR3 (N7449, N7424, N6443, N7098);
or OR4 (N7450, N7449, N5226, N5451, N359);
xor XOR2 (N7451, N7450, N5423);
or OR4 (N7452, N7445, N5214, N6719, N4867);
or OR3 (N7453, N7447, N2674, N5509);
not NOT1 (N7454, N7448);
or OR4 (N7455, N7425, N6892, N5433, N372);
buf BUF1 (N7456, N7434);
and AND3 (N7457, N7432, N14, N6812);
or OR3 (N7458, N7454, N1642, N1236);
nor NOR4 (N7459, N7451, N3770, N3706, N5099);
or OR3 (N7460, N7429, N2090, N5632);
nor NOR2 (N7461, N7460, N133);
xor XOR2 (N7462, N7458, N3002);
not NOT1 (N7463, N7440);
or OR3 (N7464, N7452, N5772, N4964);
nand NAND2 (N7465, N7464, N786);
and AND4 (N7466, N7456, N1649, N2728, N4363);
nor NOR2 (N7467, N7457, N3246);
or OR3 (N7468, N7459, N4793, N2674);
nor NOR3 (N7469, N7465, N4189, N5082);
buf BUF1 (N7470, N7461);
and AND2 (N7471, N7470, N6398);
xor XOR2 (N7472, N7462, N3650);
xor XOR2 (N7473, N7453, N6016);
nor NOR3 (N7474, N7446, N6826, N793);
not NOT1 (N7475, N7463);
nand NAND3 (N7476, N7474, N3076, N6322);
nand NAND2 (N7477, N7468, N6926);
xor XOR2 (N7478, N7471, N2081);
or OR4 (N7479, N7477, N4263, N1297, N1376);
xor XOR2 (N7480, N7469, N3753);
and AND4 (N7481, N7478, N6445, N3531, N6717);
not NOT1 (N7482, N7472);
and AND2 (N7483, N7455, N1565);
xor XOR2 (N7484, N7482, N7094);
or OR2 (N7485, N7476, N3552);
not NOT1 (N7486, N7484);
xor XOR2 (N7487, N7486, N5927);
not NOT1 (N7488, N7480);
nor NOR4 (N7489, N7475, N2063, N4514, N2492);
or OR2 (N7490, N7473, N2670);
nand NAND3 (N7491, N7483, N7162, N4324);
xor XOR2 (N7492, N7489, N7338);
or OR4 (N7493, N7492, N4056, N2590, N433);
xor XOR2 (N7494, N7487, N5795);
and AND3 (N7495, N7494, N489, N3745);
nor NOR4 (N7496, N7481, N139, N3250, N6114);
buf BUF1 (N7497, N7495);
nor NOR3 (N7498, N7493, N2625, N6933);
and AND2 (N7499, N7490, N3960);
nor NOR3 (N7500, N7497, N4939, N3762);
not NOT1 (N7501, N7499);
not NOT1 (N7502, N7500);
xor XOR2 (N7503, N7491, N1546);
and AND3 (N7504, N7467, N5721, N7245);
or OR2 (N7505, N7485, N5141);
nand NAND3 (N7506, N7496, N7460, N2762);
nand NAND2 (N7507, N7506, N1619);
or OR3 (N7508, N7479, N4259, N2821);
and AND4 (N7509, N7501, N5020, N804, N7463);
buf BUF1 (N7510, N7509);
xor XOR2 (N7511, N7498, N3274);
not NOT1 (N7512, N7508);
xor XOR2 (N7513, N7504, N5810);
xor XOR2 (N7514, N7512, N1590);
and AND3 (N7515, N7488, N4050, N2115);
nand NAND2 (N7516, N7513, N6637);
xor XOR2 (N7517, N7515, N3431);
xor XOR2 (N7518, N7507, N2482);
nor NOR4 (N7519, N7516, N7264, N2601, N4815);
nor NOR3 (N7520, N7505, N2967, N5228);
xor XOR2 (N7521, N7502, N1075);
or OR3 (N7522, N7519, N5832, N2956);
and AND2 (N7523, N7517, N559);
and AND4 (N7524, N7503, N3720, N1021, N413);
nor NOR4 (N7525, N7520, N2612, N6814, N4160);
nand NAND2 (N7526, N7522, N5653);
and AND3 (N7527, N7523, N3701, N3401);
xor XOR2 (N7528, N7524, N4625);
nand NAND2 (N7529, N7510, N6397);
nor NOR3 (N7530, N7521, N1002, N3892);
buf BUF1 (N7531, N7466);
or OR3 (N7532, N7528, N5360, N336);
buf BUF1 (N7533, N7527);
xor XOR2 (N7534, N7531, N6047);
buf BUF1 (N7535, N7511);
not NOT1 (N7536, N7529);
buf BUF1 (N7537, N7535);
nand NAND3 (N7538, N7526, N289, N6590);
xor XOR2 (N7539, N7536, N3282);
nand NAND2 (N7540, N7514, N288);
buf BUF1 (N7541, N7540);
nand NAND2 (N7542, N7518, N804);
and AND3 (N7543, N7530, N3182, N6810);
not NOT1 (N7544, N7541);
nand NAND2 (N7545, N7534, N3677);
and AND4 (N7546, N7545, N5241, N3901, N301);
and AND2 (N7547, N7532, N7072);
not NOT1 (N7548, N7533);
not NOT1 (N7549, N7525);
xor XOR2 (N7550, N7546, N1306);
or OR4 (N7551, N7537, N1061, N5392, N2026);
xor XOR2 (N7552, N7549, N6125);
or OR2 (N7553, N7544, N780);
and AND4 (N7554, N7548, N5916, N2018, N1222);
not NOT1 (N7555, N7543);
not NOT1 (N7556, N7539);
and AND2 (N7557, N7552, N2654);
buf BUF1 (N7558, N7547);
and AND2 (N7559, N7557, N912);
nand NAND4 (N7560, N7558, N1523, N6335, N5019);
not NOT1 (N7561, N7538);
not NOT1 (N7562, N7542);
xor XOR2 (N7563, N7550, N1859);
nor NOR3 (N7564, N7562, N7537, N4896);
buf BUF1 (N7565, N7560);
nor NOR4 (N7566, N7553, N58, N339, N1882);
buf BUF1 (N7567, N7554);
nor NOR4 (N7568, N7556, N1560, N5895, N3759);
nor NOR2 (N7569, N7563, N4046);
nand NAND2 (N7570, N7551, N3653);
nand NAND2 (N7571, N7567, N2097);
xor XOR2 (N7572, N7571, N3879);
and AND3 (N7573, N7561, N5287, N1385);
nand NAND2 (N7574, N7572, N4858);
or OR3 (N7575, N7564, N5573, N571);
buf BUF1 (N7576, N7566);
or OR4 (N7577, N7569, N4779, N653, N5382);
nand NAND3 (N7578, N7565, N3269, N4823);
buf BUF1 (N7579, N7577);
or OR2 (N7580, N7570, N3732);
and AND2 (N7581, N7574, N3440);
not NOT1 (N7582, N7573);
nand NAND4 (N7583, N7575, N4065, N5547, N827);
xor XOR2 (N7584, N7555, N7427);
xor XOR2 (N7585, N7580, N621);
or OR3 (N7586, N7568, N6273, N7164);
nand NAND3 (N7587, N7581, N631, N5881);
nand NAND3 (N7588, N7585, N1405, N975);
or OR2 (N7589, N7586, N60);
buf BUF1 (N7590, N7559);
buf BUF1 (N7591, N7578);
or OR2 (N7592, N7584, N2835);
or OR4 (N7593, N7591, N6777, N4949, N4804);
xor XOR2 (N7594, N7590, N2412);
nand NAND3 (N7595, N7588, N6282, N1703);
and AND3 (N7596, N7579, N7378, N6674);
xor XOR2 (N7597, N7593, N6103);
not NOT1 (N7598, N7596);
nand NAND3 (N7599, N7592, N7139, N3542);
nor NOR2 (N7600, N7594, N3546);
buf BUF1 (N7601, N7589);
xor XOR2 (N7602, N7587, N5519);
buf BUF1 (N7603, N7599);
and AND2 (N7604, N7597, N3775);
xor XOR2 (N7605, N7576, N1086);
or OR4 (N7606, N7602, N7446, N3749, N3237);
xor XOR2 (N7607, N7603, N2891);
nand NAND4 (N7608, N7582, N837, N1009, N7428);
and AND3 (N7609, N7600, N3695, N2859);
and AND4 (N7610, N7595, N2402, N69, N1651);
and AND3 (N7611, N7610, N3001, N3808);
not NOT1 (N7612, N7601);
and AND4 (N7613, N7609, N7472, N4155, N3215);
or OR2 (N7614, N7607, N150);
buf BUF1 (N7615, N7606);
buf BUF1 (N7616, N7583);
nor NOR3 (N7617, N7616, N3916, N1081);
or OR4 (N7618, N7611, N3599, N6651, N4957);
xor XOR2 (N7619, N7604, N3711);
buf BUF1 (N7620, N7612);
nor NOR2 (N7621, N7617, N6279);
buf BUF1 (N7622, N7619);
nor NOR2 (N7623, N7615, N315);
nand NAND4 (N7624, N7598, N7191, N1644, N3862);
nand NAND3 (N7625, N7614, N5429, N3911);
or OR4 (N7626, N7621, N2580, N4119, N6207);
and AND4 (N7627, N7622, N6238, N4347, N5553);
or OR2 (N7628, N7618, N265);
nand NAND4 (N7629, N7624, N2330, N800, N3402);
xor XOR2 (N7630, N7625, N4022);
and AND3 (N7631, N7623, N2049, N734);
nor NOR3 (N7632, N7605, N3438, N6594);
buf BUF1 (N7633, N7632);
buf BUF1 (N7634, N7627);
nand NAND3 (N7635, N7634, N1473, N5636);
nand NAND4 (N7636, N7613, N7569, N5005, N6582);
xor XOR2 (N7637, N7626, N7534);
nand NAND3 (N7638, N7635, N2906, N4911);
and AND4 (N7639, N7636, N3610, N6331, N4761);
and AND4 (N7640, N7629, N644, N2854, N4088);
not NOT1 (N7641, N7633);
not NOT1 (N7642, N7637);
xor XOR2 (N7643, N7642, N5219);
not NOT1 (N7644, N7631);
not NOT1 (N7645, N7638);
buf BUF1 (N7646, N7620);
or OR3 (N7647, N7646, N3034, N3105);
not NOT1 (N7648, N7628);
not NOT1 (N7649, N7639);
buf BUF1 (N7650, N7648);
nand NAND2 (N7651, N7647, N4226);
and AND4 (N7652, N7644, N951, N2499, N5081);
not NOT1 (N7653, N7630);
nor NOR2 (N7654, N7650, N24);
and AND4 (N7655, N7608, N2852, N5085, N5936);
not NOT1 (N7656, N7654);
or OR2 (N7657, N7652, N2844);
or OR3 (N7658, N7640, N1671, N3912);
and AND4 (N7659, N7649, N5269, N2738, N1044);
nor NOR3 (N7660, N7653, N4345, N53);
xor XOR2 (N7661, N7641, N2092);
buf BUF1 (N7662, N7658);
or OR4 (N7663, N7651, N2341, N1082, N38);
not NOT1 (N7664, N7645);
and AND4 (N7665, N7664, N358, N1334, N21);
nand NAND3 (N7666, N7659, N5092, N6774);
xor XOR2 (N7667, N7643, N5616);
and AND3 (N7668, N7661, N5766, N5972);
nor NOR4 (N7669, N7655, N7151, N3057, N3400);
or OR2 (N7670, N7667, N3460);
nor NOR4 (N7671, N7662, N2308, N5394, N7629);
and AND3 (N7672, N7663, N4466, N983);
buf BUF1 (N7673, N7670);
and AND4 (N7674, N7668, N7026, N7542, N1663);
nor NOR3 (N7675, N7665, N2243, N4470);
not NOT1 (N7676, N7660);
nor NOR2 (N7677, N7674, N377);
or OR3 (N7678, N7666, N7265, N1903);
buf BUF1 (N7679, N7676);
nor NOR2 (N7680, N7679, N3836);
xor XOR2 (N7681, N7678, N5993);
nor NOR2 (N7682, N7672, N530);
and AND4 (N7683, N7671, N6264, N6834, N1925);
nor NOR3 (N7684, N7681, N6888, N280);
nor NOR3 (N7685, N7673, N7170, N2835);
or OR4 (N7686, N7683, N536, N1472, N2195);
nand NAND3 (N7687, N7682, N3917, N1244);
not NOT1 (N7688, N7675);
not NOT1 (N7689, N7685);
not NOT1 (N7690, N7656);
buf BUF1 (N7691, N7686);
or OR3 (N7692, N7687, N1873, N2936);
not NOT1 (N7693, N7688);
buf BUF1 (N7694, N7691);
and AND4 (N7695, N7677, N3035, N1588, N3334);
or OR4 (N7696, N7680, N2087, N7083, N5596);
and AND4 (N7697, N7684, N1459, N2335, N7140);
nor NOR4 (N7698, N7690, N4380, N1105, N3064);
not NOT1 (N7699, N7695);
and AND3 (N7700, N7697, N780, N7028);
xor XOR2 (N7701, N7657, N4002);
not NOT1 (N7702, N7700);
not NOT1 (N7703, N7698);
nor NOR3 (N7704, N7703, N7450, N7100);
buf BUF1 (N7705, N7702);
and AND4 (N7706, N7699, N7579, N2469, N5387);
nand NAND4 (N7707, N7692, N7434, N7347, N3464);
xor XOR2 (N7708, N7689, N3919);
xor XOR2 (N7709, N7694, N7499);
buf BUF1 (N7710, N7696);
and AND4 (N7711, N7704, N3592, N1030, N6428);
nor NOR3 (N7712, N7707, N5286, N4388);
and AND4 (N7713, N7669, N5592, N3091, N6930);
xor XOR2 (N7714, N7708, N6440);
nor NOR4 (N7715, N7712, N3901, N5976, N6198);
buf BUF1 (N7716, N7705);
not NOT1 (N7717, N7715);
and AND3 (N7718, N7706, N6729, N4297);
nand NAND2 (N7719, N7709, N431);
and AND2 (N7720, N7693, N654);
xor XOR2 (N7721, N7710, N7031);
or OR3 (N7722, N7721, N3738, N6014);
buf BUF1 (N7723, N7701);
nand NAND3 (N7724, N7716, N1207, N7506);
nor NOR2 (N7725, N7714, N1565);
not NOT1 (N7726, N7720);
not NOT1 (N7727, N7724);
or OR2 (N7728, N7719, N893);
not NOT1 (N7729, N7726);
xor XOR2 (N7730, N7728, N6934);
xor XOR2 (N7731, N7713, N2655);
not NOT1 (N7732, N7731);
or OR3 (N7733, N7723, N2360, N2715);
nand NAND2 (N7734, N7727, N5425);
and AND4 (N7735, N7730, N3659, N6706, N834);
nand NAND3 (N7736, N7722, N5778, N3983);
or OR3 (N7737, N7733, N5586, N1743);
xor XOR2 (N7738, N7734, N4093);
xor XOR2 (N7739, N7732, N221);
buf BUF1 (N7740, N7735);
nand NAND2 (N7741, N7738, N6408);
and AND3 (N7742, N7736, N696, N1356);
nor NOR2 (N7743, N7717, N875);
or OR3 (N7744, N7741, N3075, N2988);
or OR3 (N7745, N7742, N3162, N4363);
nand NAND3 (N7746, N7725, N2438, N1365);
xor XOR2 (N7747, N7718, N1684);
or OR4 (N7748, N7743, N6994, N152, N2507);
xor XOR2 (N7749, N7729, N6467);
xor XOR2 (N7750, N7739, N7199);
and AND4 (N7751, N7750, N4898, N5030, N447);
nand NAND2 (N7752, N7746, N7013);
nor NOR4 (N7753, N7748, N2888, N301, N4098);
buf BUF1 (N7754, N7752);
buf BUF1 (N7755, N7747);
and AND2 (N7756, N7753, N2834);
and AND4 (N7757, N7755, N3707, N7551, N2468);
buf BUF1 (N7758, N7754);
buf BUF1 (N7759, N7711);
or OR4 (N7760, N7744, N5450, N3539, N7487);
not NOT1 (N7761, N7758);
nor NOR2 (N7762, N7756, N7271);
xor XOR2 (N7763, N7745, N4551);
and AND2 (N7764, N7740, N6673);
xor XOR2 (N7765, N7760, N279);
nand NAND4 (N7766, N7757, N4834, N2513, N1265);
not NOT1 (N7767, N7766);
nor NOR3 (N7768, N7762, N1145, N4254);
buf BUF1 (N7769, N7765);
or OR4 (N7770, N7763, N2563, N4318, N5610);
buf BUF1 (N7771, N7770);
buf BUF1 (N7772, N7769);
not NOT1 (N7773, N7767);
nand NAND3 (N7774, N7764, N4501, N508);
xor XOR2 (N7775, N7761, N600);
or OR2 (N7776, N7749, N2082);
buf BUF1 (N7777, N7759);
or OR2 (N7778, N7775, N3275);
xor XOR2 (N7779, N7778, N5457);
nand NAND4 (N7780, N7777, N6911, N2243, N4586);
or OR3 (N7781, N7776, N4979, N6918);
nand NAND4 (N7782, N7771, N877, N5083, N356);
buf BUF1 (N7783, N7781);
or OR4 (N7784, N7780, N541, N3105, N7436);
nor NOR4 (N7785, N7768, N5629, N4402, N3428);
buf BUF1 (N7786, N7751);
nand NAND2 (N7787, N7772, N4201);
not NOT1 (N7788, N7773);
nand NAND3 (N7789, N7779, N663, N4423);
and AND4 (N7790, N7785, N219, N131, N201);
or OR3 (N7791, N7788, N6378, N1729);
nand NAND2 (N7792, N7783, N7587);
nor NOR4 (N7793, N7774, N7740, N854, N2836);
not NOT1 (N7794, N7793);
not NOT1 (N7795, N7787);
nor NOR2 (N7796, N7737, N6473);
xor XOR2 (N7797, N7792, N2446);
or OR2 (N7798, N7784, N2864);
nand NAND3 (N7799, N7786, N7044, N4654);
nand NAND2 (N7800, N7797, N7505);
or OR3 (N7801, N7790, N3922, N3039);
not NOT1 (N7802, N7798);
and AND3 (N7803, N7794, N2706, N1645);
and AND2 (N7804, N7800, N6292);
xor XOR2 (N7805, N7799, N269);
nor NOR3 (N7806, N7801, N4695, N553);
buf BUF1 (N7807, N7796);
nand NAND3 (N7808, N7803, N2261, N73);
nor NOR2 (N7809, N7807, N1030);
and AND4 (N7810, N7791, N7718, N2814, N1506);
or OR4 (N7811, N7802, N5844, N3961, N411);
xor XOR2 (N7812, N7811, N2554);
xor XOR2 (N7813, N7806, N1177);
xor XOR2 (N7814, N7810, N1711);
and AND2 (N7815, N7812, N2203);
buf BUF1 (N7816, N7804);
nand NAND2 (N7817, N7782, N7046);
or OR2 (N7818, N7795, N5950);
and AND4 (N7819, N7805, N6062, N4651, N3538);
xor XOR2 (N7820, N7808, N2807);
nand NAND2 (N7821, N7789, N6473);
xor XOR2 (N7822, N7817, N7665);
and AND3 (N7823, N7820, N4718, N829);
buf BUF1 (N7824, N7814);
xor XOR2 (N7825, N7819, N6554);
nor NOR2 (N7826, N7821, N2105);
and AND3 (N7827, N7816, N3648, N5894);
buf BUF1 (N7828, N7815);
not NOT1 (N7829, N7813);
and AND4 (N7830, N7824, N142, N687, N3624);
and AND4 (N7831, N7829, N4909, N1298, N4452);
xor XOR2 (N7832, N7818, N6945);
buf BUF1 (N7833, N7827);
not NOT1 (N7834, N7825);
nand NAND4 (N7835, N7823, N1241, N3528, N4645);
nand NAND2 (N7836, N7828, N4883);
nand NAND3 (N7837, N7831, N5512, N2080);
nor NOR3 (N7838, N7830, N2096, N5927);
nor NOR2 (N7839, N7836, N1027);
nand NAND3 (N7840, N7839, N6926, N4576);
or OR4 (N7841, N7835, N4546, N1254, N6146);
xor XOR2 (N7842, N7838, N7163);
nor NOR4 (N7843, N7834, N257, N904, N677);
nor NOR3 (N7844, N7837, N7563, N6468);
and AND4 (N7845, N7842, N2478, N5410, N1192);
or OR3 (N7846, N7833, N4266, N6174);
buf BUF1 (N7847, N7832);
buf BUF1 (N7848, N7845);
buf BUF1 (N7849, N7822);
buf BUF1 (N7850, N7846);
not NOT1 (N7851, N7841);
buf BUF1 (N7852, N7844);
nor NOR3 (N7853, N7826, N6196, N2420);
and AND4 (N7854, N7852, N7477, N7470, N2348);
or OR3 (N7855, N7809, N1578, N7819);
or OR2 (N7856, N7855, N819);
and AND4 (N7857, N7843, N2743, N731, N1937);
not NOT1 (N7858, N7840);
nand NAND2 (N7859, N7850, N1282);
not NOT1 (N7860, N7851);
buf BUF1 (N7861, N7860);
nor NOR3 (N7862, N7853, N2116, N673);
nor NOR2 (N7863, N7857, N4236);
and AND3 (N7864, N7854, N7614, N1765);
or OR3 (N7865, N7861, N6544, N2155);
or OR3 (N7866, N7849, N4286, N6701);
buf BUF1 (N7867, N7864);
or OR3 (N7868, N7865, N7496, N6094);
not NOT1 (N7869, N7863);
buf BUF1 (N7870, N7848);
or OR4 (N7871, N7870, N1796, N2197, N6817);
nor NOR4 (N7872, N7858, N6846, N5842, N2176);
not NOT1 (N7873, N7867);
buf BUF1 (N7874, N7868);
nand NAND4 (N7875, N7869, N5775, N5579, N2386);
and AND2 (N7876, N7859, N7719);
nand NAND3 (N7877, N7872, N6383, N6109);
nand NAND4 (N7878, N7877, N1781, N864, N3504);
nand NAND4 (N7879, N7873, N3773, N4351, N3409);
nor NOR3 (N7880, N7874, N7646, N1241);
or OR2 (N7881, N7862, N5251);
buf BUF1 (N7882, N7847);
nand NAND2 (N7883, N7878, N6364);
xor XOR2 (N7884, N7866, N590);
nand NAND4 (N7885, N7876, N3567, N6428, N292);
not NOT1 (N7886, N7881);
nor NOR4 (N7887, N7879, N5504, N7583, N3095);
not NOT1 (N7888, N7882);
nor NOR3 (N7889, N7888, N5496, N909);
not NOT1 (N7890, N7887);
nor NOR2 (N7891, N7885, N6004);
nor NOR4 (N7892, N7890, N3385, N7020, N7132);
and AND2 (N7893, N7884, N889);
xor XOR2 (N7894, N7856, N7399);
nor NOR2 (N7895, N7891, N1318);
buf BUF1 (N7896, N7886);
or OR2 (N7897, N7894, N1395);
and AND4 (N7898, N7895, N6494, N1767, N7623);
buf BUF1 (N7899, N7897);
buf BUF1 (N7900, N7899);
and AND4 (N7901, N7896, N4586, N6385, N3651);
nor NOR4 (N7902, N7892, N5487, N903, N4722);
nand NAND4 (N7903, N7880, N1405, N6497, N2571);
nor NOR4 (N7904, N7901, N6821, N5730, N7565);
xor XOR2 (N7905, N7889, N1359);
buf BUF1 (N7906, N7898);
nand NAND2 (N7907, N7900, N3729);
and AND2 (N7908, N7903, N1320);
not NOT1 (N7909, N7875);
xor XOR2 (N7910, N7904, N5725);
not NOT1 (N7911, N7893);
xor XOR2 (N7912, N7907, N7227);
and AND2 (N7913, N7883, N879);
buf BUF1 (N7914, N7902);
xor XOR2 (N7915, N7912, N4921);
nor NOR4 (N7916, N7871, N779, N6586, N1069);
buf BUF1 (N7917, N7909);
buf BUF1 (N7918, N7914);
and AND2 (N7919, N7915, N2638);
not NOT1 (N7920, N7910);
xor XOR2 (N7921, N7908, N414);
buf BUF1 (N7922, N7906);
buf BUF1 (N7923, N7922);
nor NOR4 (N7924, N7920, N3337, N1351, N2107);
xor XOR2 (N7925, N7916, N294);
nor NOR2 (N7926, N7917, N7307);
xor XOR2 (N7927, N7925, N399);
nor NOR3 (N7928, N7923, N2731, N7452);
nand NAND2 (N7929, N7911, N119);
not NOT1 (N7930, N7913);
and AND3 (N7931, N7927, N851, N4400);
nand NAND3 (N7932, N7921, N7440, N5572);
xor XOR2 (N7933, N7926, N4627);
xor XOR2 (N7934, N7932, N7466);
buf BUF1 (N7935, N7905);
or OR4 (N7936, N7935, N1212, N3928, N386);
xor XOR2 (N7937, N7929, N87);
or OR3 (N7938, N7936, N4414, N1015);
buf BUF1 (N7939, N7937);
nand NAND3 (N7940, N7930, N7769, N1314);
not NOT1 (N7941, N7928);
xor XOR2 (N7942, N7934, N7311);
nor NOR3 (N7943, N7942, N2116, N6941);
nand NAND2 (N7944, N7931, N3416);
nand NAND2 (N7945, N7944, N777);
buf BUF1 (N7946, N7924);
and AND2 (N7947, N7945, N4589);
nand NAND3 (N7948, N7946, N2102, N3029);
and AND3 (N7949, N7939, N6366, N4360);
nor NOR4 (N7950, N7941, N7387, N5355, N6958);
not NOT1 (N7951, N7940);
nand NAND3 (N7952, N7943, N3502, N3802);
or OR2 (N7953, N7938, N5235);
not NOT1 (N7954, N7918);
or OR2 (N7955, N7948, N4352);
buf BUF1 (N7956, N7951);
xor XOR2 (N7957, N7950, N5575);
nand NAND3 (N7958, N7956, N2587, N2649);
buf BUF1 (N7959, N7933);
and AND4 (N7960, N7959, N5942, N2646, N3541);
not NOT1 (N7961, N7919);
buf BUF1 (N7962, N7953);
nand NAND4 (N7963, N7954, N7772, N1177, N3092);
or OR3 (N7964, N7960, N4650, N2524);
nor NOR2 (N7965, N7952, N4137);
buf BUF1 (N7966, N7963);
or OR2 (N7967, N7961, N6393);
or OR4 (N7968, N7967, N6037, N3390, N6473);
xor XOR2 (N7969, N7968, N1284);
buf BUF1 (N7970, N7957);
not NOT1 (N7971, N7969);
nor NOR2 (N7972, N7964, N5116);
buf BUF1 (N7973, N7955);
nand NAND4 (N7974, N7970, N3640, N1837, N6288);
and AND2 (N7975, N7966, N502);
or OR3 (N7976, N7965, N4864, N4205);
nor NOR4 (N7977, N7947, N3460, N7837, N3165);
nand NAND3 (N7978, N7975, N2734, N6634);
nor NOR3 (N7979, N7958, N260, N4037);
not NOT1 (N7980, N7976);
nand NAND2 (N7981, N7978, N5132);
xor XOR2 (N7982, N7974, N3860);
nor NOR4 (N7983, N7972, N32, N689, N5849);
and AND3 (N7984, N7981, N6059, N376);
or OR2 (N7985, N7979, N6413);
nor NOR3 (N7986, N7973, N6265, N2725);
nor NOR3 (N7987, N7985, N4273, N3429);
xor XOR2 (N7988, N7949, N7731);
not NOT1 (N7989, N7986);
or OR3 (N7990, N7980, N4492, N2971);
or OR4 (N7991, N7977, N561, N5750, N3615);
and AND3 (N7992, N7984, N758, N6054);
nand NAND4 (N7993, N7987, N4418, N2675, N5877);
and AND3 (N7994, N7988, N7294, N6789);
buf BUF1 (N7995, N7993);
buf BUF1 (N7996, N7994);
not NOT1 (N7997, N7995);
xor XOR2 (N7998, N7982, N2021);
or OR3 (N7999, N7989, N5559, N2604);
or OR2 (N8000, N7996, N5949);
nand NAND4 (N8001, N7962, N1184, N5043, N7592);
nor NOR2 (N8002, N8001, N2562);
buf BUF1 (N8003, N7999);
nand NAND4 (N8004, N7983, N7410, N4515, N365);
nor NOR2 (N8005, N7971, N346);
or OR3 (N8006, N8005, N6697, N7328);
or OR3 (N8007, N8003, N7597, N2088);
or OR4 (N8008, N7997, N5344, N2039, N3608);
nand NAND3 (N8009, N8007, N742, N7427);
xor XOR2 (N8010, N8002, N910);
nand NAND3 (N8011, N8004, N222, N2584);
or OR4 (N8012, N8010, N4956, N6742, N5694);
not NOT1 (N8013, N8008);
nor NOR2 (N8014, N8013, N307);
xor XOR2 (N8015, N7991, N5792);
or OR2 (N8016, N8009, N1992);
and AND3 (N8017, N8014, N5768, N7599);
xor XOR2 (N8018, N7990, N6687);
or OR3 (N8019, N8012, N869, N1963);
and AND2 (N8020, N8016, N1059);
xor XOR2 (N8021, N8020, N5658);
nor NOR3 (N8022, N8021, N6578, N4297);
nand NAND4 (N8023, N8022, N7044, N4254, N5782);
or OR2 (N8024, N7992, N756);
not NOT1 (N8025, N8015);
nand NAND3 (N8026, N7998, N4648, N1183);
or OR4 (N8027, N8019, N6138, N188, N1576);
buf BUF1 (N8028, N8027);
not NOT1 (N8029, N8024);
not NOT1 (N8030, N8000);
nand NAND4 (N8031, N8017, N6446, N634, N6031);
nor NOR2 (N8032, N8006, N5971);
or OR4 (N8033, N8032, N7607, N4331, N5376);
buf BUF1 (N8034, N8026);
xor XOR2 (N8035, N8025, N519);
not NOT1 (N8036, N8034);
or OR4 (N8037, N8023, N2600, N1602, N1300);
not NOT1 (N8038, N8018);
nand NAND4 (N8039, N8030, N4782, N1898, N4964);
nand NAND3 (N8040, N8028, N5661, N329);
nand NAND4 (N8041, N8031, N7506, N7916, N5672);
xor XOR2 (N8042, N8041, N5300);
and AND3 (N8043, N8039, N6582, N3663);
and AND3 (N8044, N8040, N5768, N6698);
or OR2 (N8045, N8043, N3329);
not NOT1 (N8046, N8044);
not NOT1 (N8047, N8029);
and AND4 (N8048, N8046, N4851, N2911, N1963);
or OR3 (N8049, N8033, N6193, N2035);
xor XOR2 (N8050, N8048, N6785);
and AND4 (N8051, N8047, N3156, N2856, N7705);
nor NOR2 (N8052, N8045, N492);
nor NOR4 (N8053, N8036, N4876, N3752, N3805);
buf BUF1 (N8054, N8035);
nand NAND4 (N8055, N8042, N6178, N7157, N934);
nand NAND3 (N8056, N8051, N5562, N7495);
nor NOR3 (N8057, N8049, N2086, N2411);
nor NOR2 (N8058, N8011, N1030);
or OR3 (N8059, N8038, N2544, N3006);
nand NAND2 (N8060, N8055, N5159);
not NOT1 (N8061, N8057);
not NOT1 (N8062, N8054);
not NOT1 (N8063, N8058);
and AND2 (N8064, N8056, N1824);
not NOT1 (N8065, N8052);
xor XOR2 (N8066, N8060, N3279);
xor XOR2 (N8067, N8037, N6572);
or OR3 (N8068, N8065, N918, N6755);
or OR2 (N8069, N8068, N2410);
buf BUF1 (N8070, N8062);
and AND3 (N8071, N8069, N3119, N7606);
and AND4 (N8072, N8053, N5293, N294, N3058);
nand NAND4 (N8073, N8059, N7370, N2244, N724);
xor XOR2 (N8074, N8071, N1815);
nor NOR4 (N8075, N8050, N5594, N4938, N6870);
not NOT1 (N8076, N8073);
buf BUF1 (N8077, N8072);
xor XOR2 (N8078, N8066, N5221);
buf BUF1 (N8079, N8074);
xor XOR2 (N8080, N8077, N2731);
nand NAND3 (N8081, N8080, N3980, N6608);
buf BUF1 (N8082, N8078);
and AND4 (N8083, N8079, N3119, N3945, N5077);
or OR4 (N8084, N8082, N5195, N1217, N6129);
and AND4 (N8085, N8064, N893, N3089, N6028);
xor XOR2 (N8086, N8076, N5972);
xor XOR2 (N8087, N8063, N3367);
or OR2 (N8088, N8070, N5409);
or OR2 (N8089, N8085, N6416);
buf BUF1 (N8090, N8087);
buf BUF1 (N8091, N8067);
or OR2 (N8092, N8061, N4916);
buf BUF1 (N8093, N8089);
buf BUF1 (N8094, N8088);
xor XOR2 (N8095, N8090, N7259);
and AND2 (N8096, N8083, N660);
or OR3 (N8097, N8092, N1004, N4766);
not NOT1 (N8098, N8095);
nor NOR2 (N8099, N8093, N6089);
xor XOR2 (N8100, N8075, N728);
or OR3 (N8101, N8096, N882, N3322);
nand NAND4 (N8102, N8084, N4916, N453, N7944);
nor NOR2 (N8103, N8081, N4365);
xor XOR2 (N8104, N8103, N6218);
buf BUF1 (N8105, N8094);
nor NOR2 (N8106, N8100, N3274);
not NOT1 (N8107, N8106);
buf BUF1 (N8108, N8086);
or OR3 (N8109, N8104, N1788, N3037);
xor XOR2 (N8110, N8099, N2215);
buf BUF1 (N8111, N8102);
buf BUF1 (N8112, N8109);
nor NOR4 (N8113, N8098, N4574, N6728, N2949);
xor XOR2 (N8114, N8113, N2909);
xor XOR2 (N8115, N8111, N3719);
not NOT1 (N8116, N8105);
nor NOR2 (N8117, N8115, N1486);
or OR4 (N8118, N8117, N2131, N7331, N3321);
not NOT1 (N8119, N8116);
xor XOR2 (N8120, N8091, N3624);
nand NAND3 (N8121, N8097, N1015, N7964);
buf BUF1 (N8122, N8119);
xor XOR2 (N8123, N8118, N2182);
nand NAND2 (N8124, N8101, N3819);
or OR3 (N8125, N8121, N5684, N2141);
and AND3 (N8126, N8108, N515, N5336);
nor NOR2 (N8127, N8112, N2068);
or OR4 (N8128, N8126, N4586, N5215, N3891);
not NOT1 (N8129, N8127);
buf BUF1 (N8130, N8124);
xor XOR2 (N8131, N8114, N7346);
nand NAND4 (N8132, N8130, N4379, N4801, N2340);
xor XOR2 (N8133, N8123, N7529);
not NOT1 (N8134, N8132);
or OR4 (N8135, N8120, N1355, N4488, N7451);
buf BUF1 (N8136, N8122);
xor XOR2 (N8137, N8131, N1874);
buf BUF1 (N8138, N8107);
and AND2 (N8139, N8133, N1844);
not NOT1 (N8140, N8138);
buf BUF1 (N8141, N8128);
not NOT1 (N8142, N8110);
or OR3 (N8143, N8129, N6481, N1167);
not NOT1 (N8144, N8140);
not NOT1 (N8145, N8136);
xor XOR2 (N8146, N8144, N4144);
and AND3 (N8147, N8134, N5716, N6914);
nand NAND2 (N8148, N8145, N6741);
or OR3 (N8149, N8148, N6222, N3855);
nor NOR2 (N8150, N8142, N6200);
and AND3 (N8151, N8150, N1141, N6770);
nor NOR4 (N8152, N8149, N5236, N3974, N5360);
nor NOR2 (N8153, N8137, N6947);
or OR2 (N8154, N8147, N5604);
and AND3 (N8155, N8146, N2503, N6987);
not NOT1 (N8156, N8152);
nor NOR4 (N8157, N8153, N6358, N4253, N6261);
buf BUF1 (N8158, N8143);
buf BUF1 (N8159, N8156);
and AND2 (N8160, N8125, N7764);
buf BUF1 (N8161, N8141);
not NOT1 (N8162, N8135);
xor XOR2 (N8163, N8155, N3629);
buf BUF1 (N8164, N8154);
not NOT1 (N8165, N8151);
or OR2 (N8166, N8165, N6520);
or OR3 (N8167, N8159, N7817, N3203);
nor NOR2 (N8168, N8166, N7423);
buf BUF1 (N8169, N8160);
and AND4 (N8170, N8162, N3443, N2484, N5391);
and AND4 (N8171, N8157, N7306, N2529, N2546);
xor XOR2 (N8172, N8169, N1147);
nand NAND4 (N8173, N8171, N7678, N3746, N3657);
nor NOR4 (N8174, N8173, N3376, N626, N710);
not NOT1 (N8175, N8139);
xor XOR2 (N8176, N8164, N2878);
nor NOR3 (N8177, N8168, N1147, N4138);
nor NOR3 (N8178, N8163, N4424, N3049);
nand NAND3 (N8179, N8158, N2485, N4149);
not NOT1 (N8180, N8172);
and AND2 (N8181, N8175, N6172);
not NOT1 (N8182, N8176);
or OR3 (N8183, N8161, N2011, N6331);
xor XOR2 (N8184, N8183, N770);
nor NOR3 (N8185, N8170, N4593, N1666);
and AND3 (N8186, N8182, N5685, N5072);
buf BUF1 (N8187, N8179);
not NOT1 (N8188, N8177);
nand NAND2 (N8189, N8187, N651);
xor XOR2 (N8190, N8180, N7413);
nor NOR2 (N8191, N8167, N531);
buf BUF1 (N8192, N8186);
nand NAND4 (N8193, N8192, N6082, N7891, N5459);
xor XOR2 (N8194, N8185, N3114);
not NOT1 (N8195, N8189);
buf BUF1 (N8196, N8194);
nor NOR2 (N8197, N8190, N1658);
nand NAND4 (N8198, N8174, N5677, N486, N96);
and AND2 (N8199, N8178, N6689);
not NOT1 (N8200, N8188);
nand NAND3 (N8201, N8195, N5285, N4488);
or OR2 (N8202, N8200, N4510);
buf BUF1 (N8203, N8199);
buf BUF1 (N8204, N8193);
nor NOR2 (N8205, N8198, N2741);
nand NAND3 (N8206, N8184, N8058, N750);
buf BUF1 (N8207, N8202);
buf BUF1 (N8208, N8181);
or OR3 (N8209, N8207, N5954, N2516);
and AND2 (N8210, N8208, N4780);
xor XOR2 (N8211, N8205, N5880);
nand NAND2 (N8212, N8197, N4592);
nand NAND2 (N8213, N8211, N2594);
nor NOR4 (N8214, N8210, N4206, N6781, N226);
or OR4 (N8215, N8203, N2960, N959, N4271);
nor NOR3 (N8216, N8212, N313, N2821);
buf BUF1 (N8217, N8215);
and AND2 (N8218, N8191, N7781);
buf BUF1 (N8219, N8196);
nor NOR4 (N8220, N8214, N15, N5946, N573);
or OR3 (N8221, N8216, N528, N6636);
and AND3 (N8222, N8206, N3129, N1487);
buf BUF1 (N8223, N8213);
buf BUF1 (N8224, N8209);
or OR2 (N8225, N8224, N2568);
nand NAND2 (N8226, N8221, N6493);
and AND4 (N8227, N8220, N4597, N5108, N2941);
buf BUF1 (N8228, N8218);
not NOT1 (N8229, N8227);
nor NOR3 (N8230, N8226, N6558, N3688);
not NOT1 (N8231, N8228);
buf BUF1 (N8232, N8217);
xor XOR2 (N8233, N8232, N3514);
buf BUF1 (N8234, N8222);
nor NOR2 (N8235, N8204, N1313);
nor NOR2 (N8236, N8231, N6938);
nand NAND4 (N8237, N8223, N4266, N6332, N3805);
not NOT1 (N8238, N8234);
nand NAND3 (N8239, N8201, N407, N5049);
and AND3 (N8240, N8225, N2464, N7073);
xor XOR2 (N8241, N8219, N8033);
not NOT1 (N8242, N8229);
or OR3 (N8243, N8237, N680, N1253);
xor XOR2 (N8244, N8230, N24);
xor XOR2 (N8245, N8243, N7005);
xor XOR2 (N8246, N8244, N755);
nor NOR4 (N8247, N8246, N4137, N683, N354);
not NOT1 (N8248, N8239);
not NOT1 (N8249, N8238);
nor NOR4 (N8250, N8240, N5412, N5073, N8233);
xor XOR2 (N8251, N2480, N3876);
xor XOR2 (N8252, N8235, N6268);
and AND4 (N8253, N8252, N5806, N795, N7862);
and AND2 (N8254, N8251, N3286);
not NOT1 (N8255, N8247);
nand NAND2 (N8256, N8242, N91);
buf BUF1 (N8257, N8255);
nor NOR2 (N8258, N8256, N5309);
or OR4 (N8259, N8253, N2267, N3824, N6179);
nand NAND4 (N8260, N8250, N6535, N727, N4141);
or OR3 (N8261, N8241, N2329, N1821);
or OR2 (N8262, N8248, N3573);
nand NAND4 (N8263, N8262, N6833, N8162, N490);
or OR2 (N8264, N8260, N6494);
not NOT1 (N8265, N8249);
or OR2 (N8266, N8265, N2982);
xor XOR2 (N8267, N8263, N3981);
nand NAND3 (N8268, N8254, N812, N3337);
xor XOR2 (N8269, N8261, N4035);
nor NOR4 (N8270, N8269, N2401, N4744, N2845);
nand NAND2 (N8271, N8245, N3943);
and AND4 (N8272, N8266, N3535, N1068, N7068);
nand NAND4 (N8273, N8267, N553, N6174, N7628);
buf BUF1 (N8274, N8268);
buf BUF1 (N8275, N8257);
xor XOR2 (N8276, N8275, N449);
not NOT1 (N8277, N8264);
or OR2 (N8278, N8259, N7680);
not NOT1 (N8279, N8236);
xor XOR2 (N8280, N8270, N5544);
and AND4 (N8281, N8258, N6644, N3050, N7078);
nor NOR3 (N8282, N8280, N2155, N3130);
not NOT1 (N8283, N8282);
not NOT1 (N8284, N8279);
nor NOR3 (N8285, N8284, N7641, N646);
or OR3 (N8286, N8276, N3355, N5816);
xor XOR2 (N8287, N8274, N6251);
not NOT1 (N8288, N8278);
and AND2 (N8289, N8285, N1236);
buf BUF1 (N8290, N8288);
nand NAND3 (N8291, N8281, N907, N1776);
xor XOR2 (N8292, N8272, N498);
nand NAND2 (N8293, N8273, N6758);
or OR4 (N8294, N8283, N4559, N6368, N3820);
and AND4 (N8295, N8290, N3977, N1948, N1009);
and AND3 (N8296, N8277, N2458, N4088);
buf BUF1 (N8297, N8271);
buf BUF1 (N8298, N8293);
nand NAND3 (N8299, N8287, N6284, N5113);
nor NOR4 (N8300, N8291, N7565, N3949, N747);
and AND4 (N8301, N8297, N7642, N3702, N3051);
nor NOR3 (N8302, N8294, N1400, N5374);
or OR3 (N8303, N8286, N5833, N1262);
buf BUF1 (N8304, N8298);
nand NAND2 (N8305, N8300, N1861);
nand NAND4 (N8306, N8301, N6408, N3264, N22);
and AND3 (N8307, N8306, N8306, N2851);
buf BUF1 (N8308, N8304);
not NOT1 (N8309, N8289);
xor XOR2 (N8310, N8296, N2728);
xor XOR2 (N8311, N8299, N7437);
and AND4 (N8312, N8292, N6229, N83, N5752);
buf BUF1 (N8313, N8310);
and AND4 (N8314, N8311, N4382, N562, N297);
not NOT1 (N8315, N8309);
not NOT1 (N8316, N8295);
buf BUF1 (N8317, N8314);
xor XOR2 (N8318, N8313, N7818);
and AND2 (N8319, N8315, N1323);
buf BUF1 (N8320, N8305);
not NOT1 (N8321, N8312);
buf BUF1 (N8322, N8318);
buf BUF1 (N8323, N8321);
not NOT1 (N8324, N8317);
nand NAND4 (N8325, N8307, N644, N3785, N3179);
buf BUF1 (N8326, N8323);
or OR3 (N8327, N8316, N8044, N2995);
nor NOR2 (N8328, N8302, N1158);
or OR3 (N8329, N8322, N8042, N897);
nand NAND3 (N8330, N8308, N1156, N6504);
buf BUF1 (N8331, N8328);
nand NAND2 (N8332, N8326, N3210);
xor XOR2 (N8333, N8330, N6180);
xor XOR2 (N8334, N8333, N4966);
buf BUF1 (N8335, N8327);
and AND4 (N8336, N8303, N885, N4760, N6316);
not NOT1 (N8337, N8329);
buf BUF1 (N8338, N8336);
nand NAND4 (N8339, N8332, N4519, N4922, N5064);
or OR4 (N8340, N8319, N2575, N6077, N7336);
and AND3 (N8341, N8324, N2761, N3682);
nand NAND3 (N8342, N8320, N880, N2946);
xor XOR2 (N8343, N8339, N5692);
not NOT1 (N8344, N8325);
or OR4 (N8345, N8331, N8254, N1591, N585);
nor NOR4 (N8346, N8337, N521, N7436, N3914);
xor XOR2 (N8347, N8334, N1836);
buf BUF1 (N8348, N8341);
or OR3 (N8349, N8340, N4767, N272);
not NOT1 (N8350, N8345);
and AND3 (N8351, N8347, N4757, N6379);
nor NOR3 (N8352, N8342, N5591, N3219);
buf BUF1 (N8353, N8343);
nand NAND2 (N8354, N8338, N603);
buf BUF1 (N8355, N8348);
and AND2 (N8356, N8355, N6550);
buf BUF1 (N8357, N8352);
or OR4 (N8358, N8349, N2904, N1112, N3389);
and AND3 (N8359, N8357, N1642, N2746);
buf BUF1 (N8360, N8356);
buf BUF1 (N8361, N8346);
or OR3 (N8362, N8353, N7365, N1585);
xor XOR2 (N8363, N8359, N1067);
and AND3 (N8364, N8351, N7238, N6853);
and AND3 (N8365, N8363, N4048, N1479);
not NOT1 (N8366, N8360);
and AND3 (N8367, N8344, N969, N423);
not NOT1 (N8368, N8361);
xor XOR2 (N8369, N8354, N155);
nand NAND2 (N8370, N8364, N6062);
or OR2 (N8371, N8365, N111);
buf BUF1 (N8372, N8358);
not NOT1 (N8373, N8335);
or OR4 (N8374, N8366, N6127, N4792, N5569);
and AND2 (N8375, N8369, N7082);
nand NAND3 (N8376, N8374, N99, N8076);
and AND4 (N8377, N8368, N100, N1022, N8054);
and AND3 (N8378, N8377, N3345, N1729);
and AND2 (N8379, N8362, N4845);
nand NAND4 (N8380, N8373, N871, N2073, N261);
xor XOR2 (N8381, N8378, N1783);
buf BUF1 (N8382, N8372);
nand NAND4 (N8383, N8367, N4339, N6851, N1267);
buf BUF1 (N8384, N8350);
not NOT1 (N8385, N8384);
xor XOR2 (N8386, N8371, N4963);
nor NOR3 (N8387, N8381, N5253, N634);
buf BUF1 (N8388, N8379);
nor NOR3 (N8389, N8380, N1684, N2820);
nand NAND3 (N8390, N8388, N146, N3394);
not NOT1 (N8391, N8386);
and AND2 (N8392, N8391, N5043);
or OR3 (N8393, N8376, N3560, N4987);
xor XOR2 (N8394, N8393, N746);
buf BUF1 (N8395, N8389);
buf BUF1 (N8396, N8370);
or OR4 (N8397, N8390, N6873, N5382, N5107);
and AND4 (N8398, N8382, N4556, N1667, N1907);
and AND2 (N8399, N8375, N5802);
nand NAND4 (N8400, N8383, N3893, N1319, N5075);
not NOT1 (N8401, N8385);
xor XOR2 (N8402, N8387, N5190);
and AND2 (N8403, N8398, N4081);
xor XOR2 (N8404, N8401, N269);
nor NOR4 (N8405, N8396, N425, N7350, N1454);
buf BUF1 (N8406, N8392);
and AND3 (N8407, N8406, N4566, N1213);
xor XOR2 (N8408, N8395, N6094);
nor NOR2 (N8409, N8397, N8103);
xor XOR2 (N8410, N8405, N4312);
and AND2 (N8411, N8400, N5786);
not NOT1 (N8412, N8409);
or OR4 (N8413, N8411, N2631, N3019, N6916);
and AND4 (N8414, N8399, N3077, N5923, N4332);
or OR2 (N8415, N8402, N6816);
or OR3 (N8416, N8413, N4424, N8173);
not NOT1 (N8417, N8415);
nand NAND4 (N8418, N8410, N6832, N6011, N6555);
and AND4 (N8419, N8414, N6911, N6346, N4497);
nand NAND2 (N8420, N8418, N3976);
nand NAND2 (N8421, N8419, N4218);
and AND2 (N8422, N8420, N2922);
xor XOR2 (N8423, N8422, N3405);
and AND3 (N8424, N8407, N6503, N3465);
or OR4 (N8425, N8416, N8317, N31, N4835);
or OR4 (N8426, N8408, N6251, N815, N4866);
not NOT1 (N8427, N8394);
not NOT1 (N8428, N8421);
buf BUF1 (N8429, N8426);
and AND3 (N8430, N8428, N912, N792);
xor XOR2 (N8431, N8424, N3190);
not NOT1 (N8432, N8425);
buf BUF1 (N8433, N8431);
buf BUF1 (N8434, N8417);
or OR2 (N8435, N8434, N2214);
nor NOR2 (N8436, N8423, N6094);
not NOT1 (N8437, N8403);
nand NAND4 (N8438, N8436, N4432, N3636, N7226);
nor NOR4 (N8439, N8404, N3210, N7076, N6941);
nor NOR4 (N8440, N8433, N5577, N619, N3970);
buf BUF1 (N8441, N8429);
or OR4 (N8442, N8438, N5883, N2699, N5280);
nor NOR3 (N8443, N8437, N2865, N8428);
and AND2 (N8444, N8443, N3450);
xor XOR2 (N8445, N8440, N4244);
or OR2 (N8446, N8435, N6876);
nor NOR3 (N8447, N8445, N4073, N3064);
buf BUF1 (N8448, N8444);
nor NOR2 (N8449, N8432, N5787);
or OR4 (N8450, N8427, N1512, N3466, N1098);
buf BUF1 (N8451, N8449);
not NOT1 (N8452, N8447);
xor XOR2 (N8453, N8439, N4691);
xor XOR2 (N8454, N8442, N7594);
nand NAND3 (N8455, N8446, N3089, N3752);
xor XOR2 (N8456, N8454, N476);
or OR3 (N8457, N8452, N5624, N1905);
nor NOR4 (N8458, N8441, N7574, N8143, N6007);
nor NOR2 (N8459, N8448, N917);
xor XOR2 (N8460, N8453, N2920);
or OR4 (N8461, N8460, N4341, N846, N3834);
xor XOR2 (N8462, N8458, N3133);
and AND4 (N8463, N8457, N1946, N4730, N6320);
or OR2 (N8464, N8463, N4668);
not NOT1 (N8465, N8464);
xor XOR2 (N8466, N8451, N946);
and AND4 (N8467, N8455, N4124, N6006, N8211);
buf BUF1 (N8468, N8459);
not NOT1 (N8469, N8466);
nand NAND3 (N8470, N8450, N1245, N5935);
nand NAND3 (N8471, N8467, N980, N6171);
and AND4 (N8472, N8462, N4041, N3731, N3402);
xor XOR2 (N8473, N8430, N7564);
xor XOR2 (N8474, N8472, N6250);
and AND4 (N8475, N8471, N5643, N617, N2723);
nand NAND2 (N8476, N8475, N2917);
buf BUF1 (N8477, N8469);
nand NAND4 (N8478, N8456, N7699, N1185, N785);
nand NAND4 (N8479, N8473, N6411, N703, N5511);
xor XOR2 (N8480, N8412, N879);
not NOT1 (N8481, N8476);
xor XOR2 (N8482, N8478, N175);
nand NAND3 (N8483, N8481, N484, N1063);
and AND2 (N8484, N8480, N7585);
or OR3 (N8485, N8482, N7327, N4169);
nor NOR4 (N8486, N8483, N5632, N5040, N6700);
buf BUF1 (N8487, N8474);
not NOT1 (N8488, N8477);
or OR4 (N8489, N8488, N5592, N5062, N7305);
not NOT1 (N8490, N8470);
nor NOR3 (N8491, N8487, N3802, N2075);
nand NAND3 (N8492, N8465, N4470, N1926);
not NOT1 (N8493, N8486);
not NOT1 (N8494, N8493);
or OR3 (N8495, N8479, N3266, N1210);
buf BUF1 (N8496, N8491);
not NOT1 (N8497, N8461);
and AND4 (N8498, N8489, N4322, N4718, N643);
nor NOR3 (N8499, N8495, N5021, N2115);
buf BUF1 (N8500, N8468);
or OR4 (N8501, N8497, N2284, N7957, N6750);
not NOT1 (N8502, N8501);
not NOT1 (N8503, N8496);
nor NOR4 (N8504, N8503, N625, N5444, N2849);
nand NAND2 (N8505, N8499, N4314);
not NOT1 (N8506, N8484);
not NOT1 (N8507, N8494);
xor XOR2 (N8508, N8498, N8077);
xor XOR2 (N8509, N8504, N1630);
nor NOR2 (N8510, N8509, N3726);
and AND2 (N8511, N8507, N3426);
nor NOR2 (N8512, N8506, N193);
buf BUF1 (N8513, N8510);
buf BUF1 (N8514, N8502);
not NOT1 (N8515, N8508);
nor NOR4 (N8516, N8500, N2368, N2744, N6048);
or OR3 (N8517, N8512, N5024, N3520);
nor NOR4 (N8518, N8490, N7360, N6839, N7829);
not NOT1 (N8519, N8516);
xor XOR2 (N8520, N8517, N3692);
nor NOR4 (N8521, N8519, N940, N5038, N1254);
nand NAND2 (N8522, N8492, N5125);
xor XOR2 (N8523, N8521, N4074);
nand NAND4 (N8524, N8511, N6531, N6387, N5929);
and AND2 (N8525, N8514, N2758);
xor XOR2 (N8526, N8485, N3099);
or OR2 (N8527, N8522, N6700);
not NOT1 (N8528, N8518);
nor NOR2 (N8529, N8524, N5772);
nand NAND4 (N8530, N8529, N6287, N3754, N3468);
not NOT1 (N8531, N8505);
nor NOR4 (N8532, N8513, N5314, N8484, N3168);
nor NOR3 (N8533, N8527, N3118, N6476);
and AND2 (N8534, N8515, N3232);
and AND2 (N8535, N8533, N8341);
xor XOR2 (N8536, N8526, N986);
nor NOR4 (N8537, N8530, N7455, N7147, N2679);
nor NOR4 (N8538, N8531, N1424, N2115, N4547);
xor XOR2 (N8539, N8520, N1389);
nor NOR4 (N8540, N8536, N7786, N2872, N7544);
or OR2 (N8541, N8539, N5670);
xor XOR2 (N8542, N8535, N4991);
or OR2 (N8543, N8525, N5654);
or OR3 (N8544, N8532, N151, N1880);
or OR2 (N8545, N8542, N8239);
not NOT1 (N8546, N8543);
nand NAND4 (N8547, N8528, N4510, N571, N6036);
nand NAND4 (N8548, N8537, N7389, N7754, N3521);
nand NAND4 (N8549, N8541, N345, N5322, N1130);
nand NAND3 (N8550, N8544, N838, N6977);
nand NAND2 (N8551, N8546, N5380);
buf BUF1 (N8552, N8534);
xor XOR2 (N8553, N8540, N6706);
not NOT1 (N8554, N8523);
and AND2 (N8555, N8551, N1232);
not NOT1 (N8556, N8552);
nand NAND2 (N8557, N8554, N8447);
and AND4 (N8558, N8555, N378, N2226, N5052);
or OR3 (N8559, N8550, N1539, N3881);
xor XOR2 (N8560, N8548, N137);
not NOT1 (N8561, N8557);
and AND2 (N8562, N8547, N313);
buf BUF1 (N8563, N8559);
nand NAND4 (N8564, N8538, N1305, N6257, N569);
xor XOR2 (N8565, N8561, N6851);
or OR2 (N8566, N8553, N4823);
or OR3 (N8567, N8566, N7104, N8010);
not NOT1 (N8568, N8558);
xor XOR2 (N8569, N8562, N8289);
or OR3 (N8570, N8549, N7140, N7715);
or OR3 (N8571, N8563, N928, N5283);
buf BUF1 (N8572, N8565);
nand NAND2 (N8573, N8572, N5557);
or OR4 (N8574, N8570, N6918, N6960, N569);
not NOT1 (N8575, N8556);
not NOT1 (N8576, N8545);
buf BUF1 (N8577, N8573);
buf BUF1 (N8578, N8569);
nand NAND3 (N8579, N8567, N2040, N7371);
nor NOR3 (N8580, N8577, N5109, N2456);
or OR4 (N8581, N8568, N4659, N7485, N3265);
not NOT1 (N8582, N8578);
nand NAND4 (N8583, N8580, N4697, N950, N2091);
nor NOR4 (N8584, N8583, N2569, N1262, N4430);
not NOT1 (N8585, N8575);
nand NAND4 (N8586, N8560, N992, N3660, N6108);
buf BUF1 (N8587, N8571);
buf BUF1 (N8588, N8574);
nand NAND2 (N8589, N8576, N999);
not NOT1 (N8590, N8584);
buf BUF1 (N8591, N8586);
buf BUF1 (N8592, N8589);
not NOT1 (N8593, N8590);
nor NOR3 (N8594, N8591, N7384, N3167);
not NOT1 (N8595, N8592);
buf BUF1 (N8596, N8594);
nor NOR4 (N8597, N8564, N7520, N4580, N7393);
xor XOR2 (N8598, N8582, N4469);
or OR2 (N8599, N8597, N4936);
not NOT1 (N8600, N8595);
nand NAND2 (N8601, N8593, N6846);
not NOT1 (N8602, N8601);
not NOT1 (N8603, N8585);
xor XOR2 (N8604, N8587, N6181);
and AND4 (N8605, N8599, N6280, N2258, N5579);
nand NAND3 (N8606, N8605, N5450, N1464);
nor NOR4 (N8607, N8602, N6753, N449, N5861);
nor NOR4 (N8608, N8603, N32, N6470, N6411);
or OR3 (N8609, N8600, N5911, N3456);
xor XOR2 (N8610, N8606, N7997);
not NOT1 (N8611, N8610);
or OR4 (N8612, N8581, N6100, N5681, N7865);
or OR4 (N8613, N8607, N1734, N6507, N1486);
or OR2 (N8614, N8613, N7565);
buf BUF1 (N8615, N8596);
and AND4 (N8616, N8579, N4403, N7593, N5430);
nand NAND3 (N8617, N8598, N4159, N5531);
xor XOR2 (N8618, N8614, N7528);
nor NOR3 (N8619, N8609, N1778, N7308);
buf BUF1 (N8620, N8611);
not NOT1 (N8621, N8619);
and AND4 (N8622, N8617, N5107, N363, N1540);
and AND3 (N8623, N8621, N6192, N3614);
xor XOR2 (N8624, N8623, N770);
nor NOR4 (N8625, N8604, N1128, N2494, N1737);
or OR4 (N8626, N8608, N4041, N3322, N2399);
or OR3 (N8627, N8615, N2331, N2995);
or OR2 (N8628, N8588, N7280);
xor XOR2 (N8629, N8626, N3050);
buf BUF1 (N8630, N8628);
and AND3 (N8631, N8616, N3794, N566);
nor NOR2 (N8632, N8625, N2551);
xor XOR2 (N8633, N8612, N4905);
nor NOR3 (N8634, N8633, N807, N8310);
not NOT1 (N8635, N8630);
or OR4 (N8636, N8629, N5778, N5565, N3476);
nand NAND2 (N8637, N8618, N1589);
not NOT1 (N8638, N8631);
not NOT1 (N8639, N8632);
buf BUF1 (N8640, N8637);
xor XOR2 (N8641, N8620, N5912);
or OR2 (N8642, N8640, N6357);
and AND2 (N8643, N8638, N7370);
or OR4 (N8644, N8636, N3718, N4665, N7161);
buf BUF1 (N8645, N8639);
xor XOR2 (N8646, N8627, N6487);
or OR3 (N8647, N8642, N6818, N1583);
nand NAND2 (N8648, N8635, N7045);
not NOT1 (N8649, N8647);
not NOT1 (N8650, N8641);
nand NAND3 (N8651, N8649, N6838, N882);
nand NAND3 (N8652, N8650, N7204, N2350);
nor NOR2 (N8653, N8624, N7156);
xor XOR2 (N8654, N8652, N2364);
nor NOR2 (N8655, N8653, N5887);
nand NAND3 (N8656, N8643, N3338, N7791);
not NOT1 (N8657, N8656);
xor XOR2 (N8658, N8646, N3043);
nand NAND2 (N8659, N8655, N2689);
nand NAND3 (N8660, N8657, N7328, N5652);
nand NAND4 (N8661, N8634, N3180, N7079, N2897);
or OR4 (N8662, N8651, N8433, N4038, N275);
nor NOR4 (N8663, N8645, N7363, N6538, N2656);
buf BUF1 (N8664, N8662);
xor XOR2 (N8665, N8664, N943);
nand NAND3 (N8666, N8644, N1189, N2669);
and AND4 (N8667, N8622, N1638, N5614, N5254);
nand NAND4 (N8668, N8666, N5092, N8344, N4131);
buf BUF1 (N8669, N8660);
not NOT1 (N8670, N8648);
xor XOR2 (N8671, N8668, N6582);
and AND3 (N8672, N8658, N4435, N5800);
nor NOR2 (N8673, N8665, N4760);
or OR2 (N8674, N8670, N5492);
xor XOR2 (N8675, N8667, N567);
buf BUF1 (N8676, N8672);
nand NAND3 (N8677, N8676, N1701, N5861);
nand NAND4 (N8678, N8674, N6357, N5323, N1231);
nor NOR2 (N8679, N8663, N3449);
nor NOR3 (N8680, N8669, N7177, N5115);
and AND2 (N8681, N8679, N3572);
and AND2 (N8682, N8661, N7955);
and AND2 (N8683, N8678, N4539);
xor XOR2 (N8684, N8675, N256);
xor XOR2 (N8685, N8673, N4915);
and AND2 (N8686, N8659, N2148);
and AND4 (N8687, N8671, N4150, N4016, N5647);
buf BUF1 (N8688, N8683);
buf BUF1 (N8689, N8685);
not NOT1 (N8690, N8654);
nor NOR3 (N8691, N8677, N735, N3712);
or OR3 (N8692, N8689, N2702, N2080);
and AND3 (N8693, N8680, N5132, N1320);
nand NAND3 (N8694, N8688, N5125, N4461);
or OR2 (N8695, N8691, N3829);
nand NAND2 (N8696, N8690, N2151);
buf BUF1 (N8697, N8694);
nor NOR2 (N8698, N8695, N7900);
nand NAND2 (N8699, N8698, N8248);
xor XOR2 (N8700, N8696, N8027);
or OR2 (N8701, N8686, N5913);
nand NAND2 (N8702, N8682, N531);
not NOT1 (N8703, N8681);
nand NAND4 (N8704, N8687, N517, N5650, N629);
nand NAND3 (N8705, N8699, N5073, N6832);
or OR4 (N8706, N8697, N5050, N8642, N2095);
buf BUF1 (N8707, N8700);
xor XOR2 (N8708, N8701, N2562);
xor XOR2 (N8709, N8708, N6717);
and AND3 (N8710, N8709, N4509, N3851);
nor NOR4 (N8711, N8707, N6237, N4836, N3962);
nand NAND3 (N8712, N8703, N4409, N2323);
not NOT1 (N8713, N8705);
and AND2 (N8714, N8713, N5764);
not NOT1 (N8715, N8711);
not NOT1 (N8716, N8692);
nor NOR4 (N8717, N8716, N6089, N5482, N7);
nand NAND3 (N8718, N8684, N8653, N2264);
not NOT1 (N8719, N8693);
or OR2 (N8720, N8718, N8711);
nand NAND3 (N8721, N8719, N7781, N6023);
nand NAND4 (N8722, N8715, N7896, N964, N7661);
nor NOR3 (N8723, N8706, N5808, N5597);
and AND4 (N8724, N8714, N6473, N1225, N7590);
and AND2 (N8725, N8721, N1978);
and AND3 (N8726, N8702, N3725, N5502);
or OR4 (N8727, N8717, N6792, N7768, N8082);
nor NOR2 (N8728, N8712, N4658);
not NOT1 (N8729, N8704);
buf BUF1 (N8730, N8720);
xor XOR2 (N8731, N8726, N5314);
xor XOR2 (N8732, N8723, N7271);
or OR2 (N8733, N8722, N7501);
xor XOR2 (N8734, N8710, N1168);
xor XOR2 (N8735, N8729, N3651);
and AND4 (N8736, N8727, N8101, N2312, N1702);
xor XOR2 (N8737, N8736, N8286);
buf BUF1 (N8738, N8730);
buf BUF1 (N8739, N8735);
nand NAND3 (N8740, N8739, N3663, N7478);
or OR2 (N8741, N8732, N7229);
nand NAND4 (N8742, N8733, N4261, N8448, N3243);
nand NAND4 (N8743, N8738, N3438, N920, N2164);
xor XOR2 (N8744, N8728, N1631);
xor XOR2 (N8745, N8740, N3570);
nor NOR3 (N8746, N8725, N4556, N7569);
and AND2 (N8747, N8741, N7834);
nor NOR2 (N8748, N8737, N3153);
not NOT1 (N8749, N8744);
buf BUF1 (N8750, N8749);
or OR2 (N8751, N8724, N5452);
nor NOR4 (N8752, N8746, N2560, N5090, N2618);
or OR2 (N8753, N8731, N3414);
buf BUF1 (N8754, N8750);
or OR4 (N8755, N8753, N7307, N5572, N7108);
not NOT1 (N8756, N8734);
not NOT1 (N8757, N8755);
nand NAND2 (N8758, N8754, N7001);
xor XOR2 (N8759, N8745, N1592);
nor NOR2 (N8760, N8742, N2850);
xor XOR2 (N8761, N8752, N5768);
buf BUF1 (N8762, N8760);
buf BUF1 (N8763, N8743);
buf BUF1 (N8764, N8763);
buf BUF1 (N8765, N8759);
buf BUF1 (N8766, N8757);
or OR2 (N8767, N8751, N3553);
xor XOR2 (N8768, N8765, N8590);
or OR3 (N8769, N8767, N4233, N7044);
not NOT1 (N8770, N8761);
xor XOR2 (N8771, N8747, N742);
and AND2 (N8772, N8771, N383);
or OR4 (N8773, N8766, N523, N6904, N890);
nor NOR3 (N8774, N8758, N7287, N5862);
and AND3 (N8775, N8774, N5671, N7367);
xor XOR2 (N8776, N8762, N831);
not NOT1 (N8777, N8775);
buf BUF1 (N8778, N8772);
nor NOR3 (N8779, N8773, N7155, N641);
buf BUF1 (N8780, N8777);
xor XOR2 (N8781, N8778, N7954);
not NOT1 (N8782, N8769);
xor XOR2 (N8783, N8748, N2731);
or OR3 (N8784, N8782, N8514, N3210);
nor NOR3 (N8785, N8779, N8646, N3521);
buf BUF1 (N8786, N8780);
xor XOR2 (N8787, N8756, N317);
buf BUF1 (N8788, N8764);
not NOT1 (N8789, N8768);
buf BUF1 (N8790, N8781);
xor XOR2 (N8791, N8784, N2501);
not NOT1 (N8792, N8770);
buf BUF1 (N8793, N8789);
and AND4 (N8794, N8790, N386, N2884, N8401);
or OR4 (N8795, N8793, N5876, N5950, N5407);
and AND4 (N8796, N8795, N7076, N5946, N800);
buf BUF1 (N8797, N8788);
nor NOR2 (N8798, N8783, N7054);
nand NAND4 (N8799, N8787, N7055, N5615, N5896);
nor NOR3 (N8800, N8797, N6113, N5508);
nor NOR3 (N8801, N8799, N8181, N5940);
buf BUF1 (N8802, N8786);
nand NAND3 (N8803, N8800, N7157, N7018);
buf BUF1 (N8804, N8802);
or OR4 (N8805, N8801, N4919, N1321, N6176);
and AND3 (N8806, N8792, N2634, N4889);
and AND3 (N8807, N8804, N4924, N2012);
buf BUF1 (N8808, N8794);
buf BUF1 (N8809, N8785);
not NOT1 (N8810, N8791);
xor XOR2 (N8811, N8806, N7229);
or OR3 (N8812, N8811, N8148, N7401);
xor XOR2 (N8813, N8805, N6105);
nand NAND4 (N8814, N8813, N723, N5131, N7425);
or OR2 (N8815, N8810, N1860);
nor NOR2 (N8816, N8812, N2556);
nor NOR3 (N8817, N8798, N6819, N2138);
nand NAND3 (N8818, N8809, N2476, N1736);
not NOT1 (N8819, N8796);
xor XOR2 (N8820, N8818, N6604);
nor NOR4 (N8821, N8807, N3739, N7302, N6335);
nor NOR2 (N8822, N8814, N7333);
and AND4 (N8823, N8815, N2522, N2342, N4218);
buf BUF1 (N8824, N8823);
not NOT1 (N8825, N8820);
buf BUF1 (N8826, N8816);
nand NAND3 (N8827, N8821, N4768, N540);
not NOT1 (N8828, N8824);
not NOT1 (N8829, N8817);
nand NAND4 (N8830, N8825, N3571, N3515, N2657);
nand NAND4 (N8831, N8828, N2274, N761, N906);
not NOT1 (N8832, N8827);
xor XOR2 (N8833, N8776, N7838);
buf BUF1 (N8834, N8808);
nand NAND3 (N8835, N8826, N3326, N6392);
or OR2 (N8836, N8819, N8620);
nand NAND2 (N8837, N8833, N1910);
nor NOR2 (N8838, N8835, N6825);
nand NAND3 (N8839, N8838, N1826, N7193);
and AND3 (N8840, N8831, N8564, N7306);
xor XOR2 (N8841, N8829, N1613);
and AND4 (N8842, N8830, N6926, N6331, N2649);
or OR3 (N8843, N8837, N8146, N6659);
nand NAND4 (N8844, N8822, N3937, N5971, N7096);
buf BUF1 (N8845, N8836);
buf BUF1 (N8846, N8803);
nor NOR3 (N8847, N8832, N2355, N5397);
not NOT1 (N8848, N8843);
buf BUF1 (N8849, N8842);
nor NOR3 (N8850, N8840, N4913, N814);
xor XOR2 (N8851, N8845, N4964);
nand NAND4 (N8852, N8847, N5857, N5077, N4417);
and AND2 (N8853, N8846, N1145);
xor XOR2 (N8854, N8851, N180);
xor XOR2 (N8855, N8848, N7162);
nand NAND4 (N8856, N8834, N7658, N1357, N3430);
nand NAND4 (N8857, N8850, N6332, N3569, N7564);
and AND4 (N8858, N8857, N403, N7940, N7640);
nand NAND2 (N8859, N8855, N8473);
or OR2 (N8860, N8854, N7231);
nor NOR2 (N8861, N8859, N7782);
not NOT1 (N8862, N8853);
nor NOR3 (N8863, N8852, N26, N2528);
and AND2 (N8864, N8839, N1988);
nor NOR4 (N8865, N8858, N6059, N1397, N2763);
buf BUF1 (N8866, N8849);
not NOT1 (N8867, N8841);
or OR3 (N8868, N8865, N798, N1573);
nor NOR3 (N8869, N8861, N8731, N6399);
xor XOR2 (N8870, N8863, N1873);
or OR4 (N8871, N8856, N2210, N1074, N2874);
or OR2 (N8872, N8870, N4884);
or OR3 (N8873, N8868, N1232, N4000);
buf BUF1 (N8874, N8871);
and AND4 (N8875, N8869, N1048, N859, N6966);
nand NAND2 (N8876, N8872, N7536);
xor XOR2 (N8877, N8860, N6448);
xor XOR2 (N8878, N8844, N4915);
xor XOR2 (N8879, N8877, N5618);
buf BUF1 (N8880, N8867);
xor XOR2 (N8881, N8862, N2975);
nor NOR3 (N8882, N8864, N1614, N8554);
xor XOR2 (N8883, N8866, N3141);
xor XOR2 (N8884, N8883, N8677);
nor NOR2 (N8885, N8874, N5830);
and AND4 (N8886, N8878, N1909, N7041, N4626);
nor NOR4 (N8887, N8876, N4833, N5110, N1695);
nor NOR4 (N8888, N8881, N5742, N4413, N4778);
nor NOR3 (N8889, N8888, N8534, N7700);
buf BUF1 (N8890, N8875);
buf BUF1 (N8891, N8882);
xor XOR2 (N8892, N8885, N8525);
or OR2 (N8893, N8884, N5298);
and AND3 (N8894, N8880, N5153, N3792);
or OR3 (N8895, N8893, N8745, N6883);
xor XOR2 (N8896, N8891, N3304);
xor XOR2 (N8897, N8892, N1312);
nor NOR4 (N8898, N8886, N2084, N4398, N1309);
and AND4 (N8899, N8889, N4266, N7598, N7029);
buf BUF1 (N8900, N8897);
nor NOR3 (N8901, N8894, N627, N8008);
not NOT1 (N8902, N8887);
not NOT1 (N8903, N8899);
nor NOR4 (N8904, N8895, N6007, N7403, N2055);
not NOT1 (N8905, N8903);
nor NOR4 (N8906, N8898, N6377, N3689, N2306);
and AND4 (N8907, N8905, N7554, N8642, N618);
nand NAND3 (N8908, N8873, N8721, N7660);
xor XOR2 (N8909, N8907, N1099);
nand NAND3 (N8910, N8879, N2033, N890);
and AND4 (N8911, N8910, N346, N4624, N7976);
not NOT1 (N8912, N8906);
nor NOR2 (N8913, N8902, N8317);
nor NOR2 (N8914, N8912, N7090);
nor NOR3 (N8915, N8896, N1249, N4948);
xor XOR2 (N8916, N8904, N1700);
nand NAND4 (N8917, N8913, N788, N1704, N8434);
nand NAND4 (N8918, N8909, N3635, N6697, N4822);
nor NOR2 (N8919, N8918, N7017);
or OR2 (N8920, N8900, N6263);
and AND2 (N8921, N8915, N8885);
or OR3 (N8922, N8919, N5513, N332);
buf BUF1 (N8923, N8916);
buf BUF1 (N8924, N8890);
buf BUF1 (N8925, N8921);
buf BUF1 (N8926, N8917);
not NOT1 (N8927, N8922);
not NOT1 (N8928, N8926);
xor XOR2 (N8929, N8925, N2978);
buf BUF1 (N8930, N8914);
nor NOR4 (N8931, N8920, N2203, N5771, N2377);
nand NAND4 (N8932, N8923, N5302, N7756, N3291);
and AND2 (N8933, N8908, N8156);
not NOT1 (N8934, N8928);
xor XOR2 (N8935, N8930, N4819);
buf BUF1 (N8936, N8901);
nand NAND3 (N8937, N8927, N7898, N7788);
xor XOR2 (N8938, N8911, N7502);
and AND2 (N8939, N8931, N7555);
and AND3 (N8940, N8924, N3927, N3104);
buf BUF1 (N8941, N8939);
nand NAND4 (N8942, N8934, N2700, N3099, N6384);
not NOT1 (N8943, N8942);
nand NAND3 (N8944, N8936, N7619, N1199);
not NOT1 (N8945, N8932);
not NOT1 (N8946, N8944);
not NOT1 (N8947, N8945);
nand NAND3 (N8948, N8933, N607, N4621);
and AND4 (N8949, N8935, N6050, N3184, N3123);
nand NAND3 (N8950, N8929, N7768, N325);
xor XOR2 (N8951, N8946, N5611);
not NOT1 (N8952, N8940);
nand NAND2 (N8953, N8951, N98);
nor NOR3 (N8954, N8938, N3097, N1782);
and AND4 (N8955, N8937, N583, N7026, N2979);
or OR4 (N8956, N8943, N7490, N2885, N5862);
not NOT1 (N8957, N8956);
nand NAND3 (N8958, N8952, N6319, N5293);
buf BUF1 (N8959, N8950);
and AND3 (N8960, N8948, N1651, N2658);
not NOT1 (N8961, N8960);
xor XOR2 (N8962, N8959, N1701);
buf BUF1 (N8963, N8953);
or OR4 (N8964, N8962, N2735, N1121, N6819);
nand NAND2 (N8965, N8947, N2546);
or OR2 (N8966, N8949, N8737);
xor XOR2 (N8967, N8961, N4956);
or OR2 (N8968, N8941, N6888);
xor XOR2 (N8969, N8957, N7861);
xor XOR2 (N8970, N8966, N4296);
and AND2 (N8971, N8967, N931);
buf BUF1 (N8972, N8969);
nand NAND4 (N8973, N8958, N7147, N7110, N2630);
xor XOR2 (N8974, N8955, N2170);
xor XOR2 (N8975, N8964, N1951);
or OR3 (N8976, N8954, N7459, N8831);
nor NOR4 (N8977, N8968, N2766, N6010, N3099);
not NOT1 (N8978, N8970);
nor NOR4 (N8979, N8978, N3317, N4997, N5767);
nor NOR2 (N8980, N8977, N5359);
not NOT1 (N8981, N8963);
xor XOR2 (N8982, N8975, N1647);
and AND3 (N8983, N8981, N8523, N4186);
buf BUF1 (N8984, N8983);
buf BUF1 (N8985, N8971);
or OR3 (N8986, N8985, N8833, N4272);
and AND3 (N8987, N8980, N7274, N7750);
buf BUF1 (N8988, N8987);
not NOT1 (N8989, N8982);
buf BUF1 (N8990, N8973);
xor XOR2 (N8991, N8972, N4005);
nand NAND4 (N8992, N8986, N3252, N7564, N7639);
nand NAND4 (N8993, N8988, N6541, N8976, N2348);
or OR4 (N8994, N7195, N5281, N72, N2319);
xor XOR2 (N8995, N8965, N6654);
nand NAND3 (N8996, N8974, N1911, N2794);
xor XOR2 (N8997, N8984, N5432);
nor NOR2 (N8998, N8995, N6040);
xor XOR2 (N8999, N8996, N6682);
not NOT1 (N9000, N8991);
nor NOR2 (N9001, N8993, N3806);
not NOT1 (N9002, N9000);
buf BUF1 (N9003, N8998);
or OR3 (N9004, N8999, N8392, N1369);
nand NAND3 (N9005, N8994, N1767, N4451);
or OR3 (N9006, N8992, N7229, N4018);
buf BUF1 (N9007, N8979);
buf BUF1 (N9008, N9003);
nor NOR2 (N9009, N9008, N822);
nor NOR4 (N9010, N8997, N134, N8482, N7264);
nor NOR2 (N9011, N9006, N1759);
or OR2 (N9012, N8990, N8143);
xor XOR2 (N9013, N9005, N5861);
and AND3 (N9014, N9002, N5470, N2250);
not NOT1 (N9015, N9009);
xor XOR2 (N9016, N9004, N8197);
nand NAND2 (N9017, N9016, N8973);
nand NAND3 (N9018, N9012, N6318, N8663);
nand NAND4 (N9019, N9014, N2518, N1590, N5325);
buf BUF1 (N9020, N9017);
or OR4 (N9021, N9020, N7973, N50, N5042);
and AND2 (N9022, N9021, N1663);
not NOT1 (N9023, N9018);
buf BUF1 (N9024, N9015);
nand NAND3 (N9025, N9001, N8154, N6823);
not NOT1 (N9026, N9019);
not NOT1 (N9027, N9022);
nor NOR4 (N9028, N9011, N379, N5704, N6721);
and AND4 (N9029, N9010, N1845, N8306, N1650);
xor XOR2 (N9030, N9024, N5722);
or OR3 (N9031, N9007, N1079, N6471);
and AND4 (N9032, N9013, N1643, N3267, N3132);
nor NOR2 (N9033, N9023, N5010);
and AND2 (N9034, N9029, N7072);
buf BUF1 (N9035, N9033);
and AND2 (N9036, N9030, N3936);
xor XOR2 (N9037, N9025, N5967);
xor XOR2 (N9038, N9028, N2536);
xor XOR2 (N9039, N9026, N8908);
nor NOR2 (N9040, N9027, N1727);
nand NAND3 (N9041, N9035, N6916, N8120);
buf BUF1 (N9042, N8989);
nand NAND2 (N9043, N9037, N4429);
buf BUF1 (N9044, N9039);
nand NAND3 (N9045, N9036, N6439, N7795);
or OR4 (N9046, N9040, N820, N5735, N3922);
and AND4 (N9047, N9042, N8685, N4575, N2374);
xor XOR2 (N9048, N9032, N2593);
nor NOR2 (N9049, N9048, N6538);
nand NAND4 (N9050, N9041, N3665, N4242, N5979);
not NOT1 (N9051, N9034);
not NOT1 (N9052, N9031);
or OR4 (N9053, N9046, N55, N3101, N3247);
xor XOR2 (N9054, N9050, N2849);
xor XOR2 (N9055, N9043, N1968);
not NOT1 (N9056, N9052);
nor NOR4 (N9057, N9049, N6543, N8359, N836);
xor XOR2 (N9058, N9045, N7229);
xor XOR2 (N9059, N9044, N6313);
nand NAND4 (N9060, N9056, N8884, N1904, N6515);
xor XOR2 (N9061, N9054, N6571);
nand NAND3 (N9062, N9061, N5245, N6374);
nand NAND4 (N9063, N9047, N4109, N7624, N7796);
or OR2 (N9064, N9051, N6478);
buf BUF1 (N9065, N9064);
and AND3 (N9066, N9057, N8579, N9026);
xor XOR2 (N9067, N9060, N9028);
xor XOR2 (N9068, N9066, N7137);
buf BUF1 (N9069, N9065);
or OR4 (N9070, N9062, N6837, N8523, N3365);
buf BUF1 (N9071, N9070);
nand NAND3 (N9072, N9058, N1571, N3357);
or OR3 (N9073, N9063, N6055, N8177);
xor XOR2 (N9074, N9053, N9071);
xor XOR2 (N9075, N8028, N4116);
xor XOR2 (N9076, N9074, N1833);
nand NAND3 (N9077, N9068, N4178, N2116);
xor XOR2 (N9078, N9038, N8113);
not NOT1 (N9079, N9073);
nor NOR3 (N9080, N9072, N6569, N5610);
not NOT1 (N9081, N9080);
nand NAND4 (N9082, N9076, N1352, N7924, N6886);
buf BUF1 (N9083, N9082);
and AND3 (N9084, N9077, N7943, N1137);
not NOT1 (N9085, N9067);
xor XOR2 (N9086, N9079, N4506);
nor NOR2 (N9087, N9086, N3279);
nor NOR3 (N9088, N9069, N8054, N4515);
or OR4 (N9089, N9087, N9076, N3654, N1105);
or OR4 (N9090, N9055, N8415, N2147, N638);
xor XOR2 (N9091, N9085, N7803);
or OR3 (N9092, N9075, N2032, N531);
and AND4 (N9093, N9078, N8415, N3040, N6418);
xor XOR2 (N9094, N9092, N11);
and AND3 (N9095, N9059, N745, N2674);
nor NOR4 (N9096, N9093, N8888, N5922, N3020);
nor NOR4 (N9097, N9094, N3399, N1821, N7930);
nor NOR4 (N9098, N9095, N8955, N8625, N2556);
nor NOR3 (N9099, N9096, N1831, N5006);
nand NAND4 (N9100, N9090, N7920, N2902, N5286);
nor NOR2 (N9101, N9081, N3495);
buf BUF1 (N9102, N9091);
nor NOR3 (N9103, N9099, N3711, N4093);
buf BUF1 (N9104, N9098);
buf BUF1 (N9105, N9100);
nand NAND3 (N9106, N9102, N2737, N7024);
not NOT1 (N9107, N9083);
buf BUF1 (N9108, N9084);
not NOT1 (N9109, N9101);
nand NAND4 (N9110, N9109, N3157, N2036, N7001);
or OR2 (N9111, N9088, N3931);
nand NAND2 (N9112, N9111, N1826);
buf BUF1 (N9113, N9108);
not NOT1 (N9114, N9110);
not NOT1 (N9115, N9097);
xor XOR2 (N9116, N9103, N8448);
nor NOR4 (N9117, N9114, N2112, N170, N1452);
not NOT1 (N9118, N9105);
or OR4 (N9119, N9115, N7471, N473, N7731);
or OR2 (N9120, N9116, N3475);
nor NOR3 (N9121, N9117, N6021, N2384);
nand NAND2 (N9122, N9120, N8431);
buf BUF1 (N9123, N9118);
buf BUF1 (N9124, N9123);
and AND2 (N9125, N9124, N1780);
nand NAND4 (N9126, N9125, N2327, N1188, N3556);
not NOT1 (N9127, N9112);
not NOT1 (N9128, N9089);
nand NAND4 (N9129, N9119, N6322, N3289, N5549);
or OR2 (N9130, N9107, N7161);
buf BUF1 (N9131, N9121);
xor XOR2 (N9132, N9122, N2179);
buf BUF1 (N9133, N9113);
not NOT1 (N9134, N9132);
nor NOR3 (N9135, N9129, N8119, N5094);
nor NOR3 (N9136, N9133, N1479, N4076);
nor NOR3 (N9137, N9136, N7031, N114);
not NOT1 (N9138, N9135);
not NOT1 (N9139, N9134);
buf BUF1 (N9140, N9138);
not NOT1 (N9141, N9106);
nand NAND3 (N9142, N9126, N5353, N8324);
nor NOR2 (N9143, N9128, N5401);
xor XOR2 (N9144, N9139, N668);
buf BUF1 (N9145, N9127);
not NOT1 (N9146, N9104);
or OR3 (N9147, N9137, N6417, N3242);
not NOT1 (N9148, N9140);
not NOT1 (N9149, N9146);
xor XOR2 (N9150, N9145, N1167);
not NOT1 (N9151, N9150);
nand NAND3 (N9152, N9143, N6170, N3669);
not NOT1 (N9153, N9130);
or OR4 (N9154, N9144, N6364, N6346, N71);
nand NAND3 (N9155, N9154, N4528, N6520);
not NOT1 (N9156, N9131);
buf BUF1 (N9157, N9156);
nand NAND2 (N9158, N9151, N335);
and AND4 (N9159, N9142, N1152, N9031, N8672);
and AND4 (N9160, N9141, N8990, N7514, N8363);
xor XOR2 (N9161, N9158, N8568);
xor XOR2 (N9162, N9147, N1601);
buf BUF1 (N9163, N9159);
or OR2 (N9164, N9155, N5497);
not NOT1 (N9165, N9148);
buf BUF1 (N9166, N9165);
xor XOR2 (N9167, N9152, N1162);
and AND2 (N9168, N9166, N1545);
nor NOR4 (N9169, N9168, N8891, N3557, N8719);
xor XOR2 (N9170, N9149, N1440);
nand NAND4 (N9171, N9164, N7928, N8894, N1803);
xor XOR2 (N9172, N9169, N7273);
and AND2 (N9173, N9160, N6701);
buf BUF1 (N9174, N9153);
xor XOR2 (N9175, N9172, N570);
nor NOR3 (N9176, N9170, N2243, N4967);
xor XOR2 (N9177, N9163, N2746);
nand NAND3 (N9178, N9175, N7991, N7360);
not NOT1 (N9179, N9161);
nand NAND3 (N9180, N9178, N4355, N3784);
nand NAND4 (N9181, N9180, N1807, N4929, N4796);
buf BUF1 (N9182, N9174);
buf BUF1 (N9183, N9177);
not NOT1 (N9184, N9183);
and AND4 (N9185, N9157, N8316, N7892, N4938);
or OR3 (N9186, N9167, N6932, N4138);
xor XOR2 (N9187, N9186, N8111);
buf BUF1 (N9188, N9171);
and AND3 (N9189, N9162, N6922, N990);
nand NAND4 (N9190, N9179, N8603, N2362, N4325);
nand NAND3 (N9191, N9190, N3577, N8819);
not NOT1 (N9192, N9188);
and AND2 (N9193, N9191, N3103);
nor NOR2 (N9194, N9185, N5361);
buf BUF1 (N9195, N9182);
or OR3 (N9196, N9189, N3016, N7555);
xor XOR2 (N9197, N9173, N8530);
or OR3 (N9198, N9187, N7514, N406);
and AND4 (N9199, N9176, N679, N4963, N6284);
or OR4 (N9200, N9195, N4407, N2020, N1883);
xor XOR2 (N9201, N9194, N3942);
nand NAND3 (N9202, N9193, N5138, N34);
or OR3 (N9203, N9201, N30, N3592);
buf BUF1 (N9204, N9192);
nor NOR3 (N9205, N9203, N6824, N7625);
nand NAND3 (N9206, N9200, N3813, N8519);
and AND2 (N9207, N9205, N4030);
xor XOR2 (N9208, N9204, N919);
not NOT1 (N9209, N9207);
and AND4 (N9210, N9209, N1868, N1998, N3473);
xor XOR2 (N9211, N9196, N2904);
not NOT1 (N9212, N9202);
nand NAND2 (N9213, N9198, N4141);
nand NAND3 (N9214, N9208, N8148, N3206);
buf BUF1 (N9215, N9206);
buf BUF1 (N9216, N9181);
and AND3 (N9217, N9211, N7439, N4613);
nor NOR2 (N9218, N9217, N5832);
or OR2 (N9219, N9199, N4599);
buf BUF1 (N9220, N9215);
xor XOR2 (N9221, N9218, N8710);
nor NOR4 (N9222, N9212, N6675, N5763, N7864);
or OR3 (N9223, N9222, N8898, N1345);
or OR3 (N9224, N9223, N2127, N4114);
and AND4 (N9225, N9184, N6622, N1388, N5717);
xor XOR2 (N9226, N9210, N2855);
nor NOR4 (N9227, N9219, N8290, N808, N3657);
nor NOR4 (N9228, N9227, N299, N2052, N422);
nand NAND2 (N9229, N9221, N6324);
or OR3 (N9230, N9197, N4766, N4304);
xor XOR2 (N9231, N9216, N1160);
and AND3 (N9232, N9224, N355, N3288);
nand NAND2 (N9233, N9220, N6457);
or OR3 (N9234, N9213, N878, N4385);
and AND2 (N9235, N9232, N2561);
buf BUF1 (N9236, N9214);
nand NAND4 (N9237, N9236, N7547, N3583, N3428);
and AND4 (N9238, N9229, N1742, N3308, N3497);
not NOT1 (N9239, N9231);
not NOT1 (N9240, N9234);
buf BUF1 (N9241, N9230);
and AND3 (N9242, N9233, N1414, N2915);
not NOT1 (N9243, N9225);
buf BUF1 (N9244, N9226);
and AND3 (N9245, N9228, N3107, N6969);
nand NAND2 (N9246, N9245, N4774);
xor XOR2 (N9247, N9235, N5628);
not NOT1 (N9248, N9242);
nand NAND2 (N9249, N9240, N1780);
nor NOR2 (N9250, N9247, N3328);
nor NOR3 (N9251, N9237, N1434, N4058);
and AND4 (N9252, N9243, N3764, N8249, N5792);
nor NOR2 (N9253, N9250, N4726);
buf BUF1 (N9254, N9253);
or OR3 (N9255, N9254, N8451, N2758);
not NOT1 (N9256, N9246);
nor NOR4 (N9257, N9249, N8647, N8332, N5525);
not NOT1 (N9258, N9248);
buf BUF1 (N9259, N9252);
xor XOR2 (N9260, N9256, N6874);
buf BUF1 (N9261, N9258);
nand NAND4 (N9262, N9238, N6371, N5913, N295);
buf BUF1 (N9263, N9257);
and AND3 (N9264, N9244, N7492, N6822);
and AND4 (N9265, N9259, N3026, N457, N5969);
or OR3 (N9266, N9261, N5565, N6704);
or OR4 (N9267, N9265, N5405, N5803, N7763);
nand NAND2 (N9268, N9241, N8579);
buf BUF1 (N9269, N9262);
buf BUF1 (N9270, N9255);
or OR2 (N9271, N9251, N9057);
buf BUF1 (N9272, N9267);
xor XOR2 (N9273, N9271, N7500);
nand NAND4 (N9274, N9273, N2062, N5502, N3953);
xor XOR2 (N9275, N9260, N6429);
not NOT1 (N9276, N9270);
not NOT1 (N9277, N9264);
nor NOR2 (N9278, N9263, N7623);
nor NOR4 (N9279, N9269, N1437, N1777, N6818);
not NOT1 (N9280, N9275);
buf BUF1 (N9281, N9268);
and AND3 (N9282, N9278, N3964, N3691);
and AND2 (N9283, N9272, N4128);
and AND2 (N9284, N9274, N525);
buf BUF1 (N9285, N9281);
nand NAND4 (N9286, N9266, N1561, N2234, N6228);
not NOT1 (N9287, N9285);
buf BUF1 (N9288, N9277);
or OR2 (N9289, N9280, N3095);
not NOT1 (N9290, N9286);
xor XOR2 (N9291, N9287, N2549);
nand NAND4 (N9292, N9290, N6900, N249, N2356);
buf BUF1 (N9293, N9283);
and AND3 (N9294, N9293, N6724, N2467);
and AND2 (N9295, N9289, N6771);
nand NAND3 (N9296, N9292, N1818, N3945);
and AND4 (N9297, N9288, N7049, N7659, N5482);
nor NOR4 (N9298, N9291, N6120, N8865, N1844);
nor NOR3 (N9299, N9239, N718, N3761);
xor XOR2 (N9300, N9276, N4419);
not NOT1 (N9301, N9300);
nand NAND4 (N9302, N9279, N88, N3288, N1727);
buf BUF1 (N9303, N9284);
buf BUF1 (N9304, N9298);
not NOT1 (N9305, N9297);
nand NAND4 (N9306, N9301, N8067, N919, N4038);
buf BUF1 (N9307, N9294);
xor XOR2 (N9308, N9282, N4464);
or OR2 (N9309, N9308, N1352);
nor NOR4 (N9310, N9309, N5925, N2702, N8512);
buf BUF1 (N9311, N9296);
not NOT1 (N9312, N9303);
nand NAND3 (N9313, N9299, N7373, N8932);
not NOT1 (N9314, N9307);
xor XOR2 (N9315, N9311, N3024);
buf BUF1 (N9316, N9315);
buf BUF1 (N9317, N9306);
nor NOR2 (N9318, N9310, N1534);
and AND3 (N9319, N9305, N4892, N4922);
and AND2 (N9320, N9316, N5632);
buf BUF1 (N9321, N9319);
not NOT1 (N9322, N9304);
nor NOR2 (N9323, N9295, N7177);
nand NAND4 (N9324, N9314, N2072, N3716, N1231);
nor NOR3 (N9325, N9324, N4270, N7724);
xor XOR2 (N9326, N9320, N8141);
buf BUF1 (N9327, N9313);
nand NAND4 (N9328, N9318, N1133, N2898, N4867);
and AND2 (N9329, N9312, N2770);
nand NAND3 (N9330, N9328, N245, N455);
nor NOR4 (N9331, N9322, N1044, N6457, N6583);
and AND2 (N9332, N9321, N6412);
buf BUF1 (N9333, N9302);
or OR3 (N9334, N9326, N8795, N5076);
or OR4 (N9335, N9331, N7846, N532, N8981);
or OR2 (N9336, N9332, N1114);
nand NAND3 (N9337, N9329, N6422, N4528);
xor XOR2 (N9338, N9335, N3365);
and AND2 (N9339, N9323, N7490);
nand NAND4 (N9340, N9336, N8104, N4116, N215);
xor XOR2 (N9341, N9330, N4763);
and AND2 (N9342, N9339, N2476);
nor NOR4 (N9343, N9337, N3308, N5749, N3019);
xor XOR2 (N9344, N9317, N8183);
buf BUF1 (N9345, N9343);
buf BUF1 (N9346, N9333);
buf BUF1 (N9347, N9341);
or OR4 (N9348, N9340, N7846, N480, N3123);
xor XOR2 (N9349, N9348, N5392);
or OR4 (N9350, N9346, N4969, N2838, N9348);
nand NAND3 (N9351, N9344, N1913, N3661);
nor NOR2 (N9352, N9325, N6259);
or OR2 (N9353, N9342, N3157);
not NOT1 (N9354, N9338);
buf BUF1 (N9355, N9353);
nor NOR3 (N9356, N9334, N400, N9039);
xor XOR2 (N9357, N9356, N5785);
and AND4 (N9358, N9357, N1645, N5269, N7178);
and AND2 (N9359, N9345, N188);
buf BUF1 (N9360, N9354);
not NOT1 (N9361, N9327);
nor NOR3 (N9362, N9352, N1907, N9342);
nor NOR4 (N9363, N9361, N7228, N4212, N4999);
buf BUF1 (N9364, N9350);
nand NAND4 (N9365, N9364, N6843, N4087, N5987);
or OR4 (N9366, N9363, N4653, N1404, N7842);
and AND4 (N9367, N9365, N6333, N6242, N3973);
xor XOR2 (N9368, N9359, N5337);
nor NOR3 (N9369, N9367, N4296, N1184);
nand NAND3 (N9370, N9368, N1871, N5753);
buf BUF1 (N9371, N9360);
or OR4 (N9372, N9371, N4923, N4415, N1787);
not NOT1 (N9373, N9355);
and AND4 (N9374, N9372, N274, N3298, N4827);
not NOT1 (N9375, N9351);
not NOT1 (N9376, N9347);
nand NAND2 (N9377, N9375, N6035);
buf BUF1 (N9378, N9377);
buf BUF1 (N9379, N9349);
nor NOR2 (N9380, N9358, N7494);
or OR2 (N9381, N9369, N7036);
not NOT1 (N9382, N9380);
not NOT1 (N9383, N9373);
not NOT1 (N9384, N9378);
and AND2 (N9385, N9383, N6042);
nand NAND3 (N9386, N9370, N6725, N1211);
not NOT1 (N9387, N9385);
buf BUF1 (N9388, N9386);
xor XOR2 (N9389, N9388, N5121);
xor XOR2 (N9390, N9376, N5296);
and AND3 (N9391, N9382, N5861, N8037);
xor XOR2 (N9392, N9366, N2816);
and AND2 (N9393, N9392, N2839);
nand NAND2 (N9394, N9381, N8136);
buf BUF1 (N9395, N9379);
not NOT1 (N9396, N9389);
and AND3 (N9397, N9396, N7133, N5329);
buf BUF1 (N9398, N9394);
not NOT1 (N9399, N9397);
buf BUF1 (N9400, N9395);
not NOT1 (N9401, N9398);
and AND4 (N9402, N9399, N4260, N40, N639);
or OR2 (N9403, N9390, N3332);
not NOT1 (N9404, N9387);
xor XOR2 (N9405, N9403, N4931);
buf BUF1 (N9406, N9384);
or OR2 (N9407, N9401, N1706);
or OR3 (N9408, N9402, N5748, N237);
and AND2 (N9409, N9405, N8220);
xor XOR2 (N9410, N9407, N7994);
xor XOR2 (N9411, N9404, N4263);
nand NAND3 (N9412, N9410, N8503, N8123);
buf BUF1 (N9413, N9412);
nor NOR3 (N9414, N9400, N8112, N4343);
buf BUF1 (N9415, N9409);
not NOT1 (N9416, N9415);
or OR3 (N9417, N9374, N6350, N4251);
xor XOR2 (N9418, N9391, N3145);
or OR2 (N9419, N9408, N2993);
and AND3 (N9420, N9419, N9277, N3180);
and AND2 (N9421, N9416, N5567);
xor XOR2 (N9422, N9414, N1816);
xor XOR2 (N9423, N9418, N3499);
nor NOR2 (N9424, N9423, N9074);
xor XOR2 (N9425, N9406, N918);
xor XOR2 (N9426, N9425, N5553);
or OR4 (N9427, N9420, N8290, N6515, N7260);
xor XOR2 (N9428, N9411, N211);
and AND3 (N9429, N9421, N3723, N5145);
nor NOR4 (N9430, N9426, N6715, N8733, N4792);
buf BUF1 (N9431, N9424);
nor NOR2 (N9432, N9428, N7235);
and AND4 (N9433, N9422, N7317, N804, N5161);
nand NAND3 (N9434, N9417, N3487, N4947);
buf BUF1 (N9435, N9362);
buf BUF1 (N9436, N9413);
nand NAND3 (N9437, N9393, N8998, N4957);
nor NOR3 (N9438, N9427, N842, N8108);
or OR3 (N9439, N9436, N4104, N1592);
nor NOR2 (N9440, N9429, N1401);
or OR3 (N9441, N9439, N2171, N517);
or OR2 (N9442, N9430, N6703);
not NOT1 (N9443, N9433);
and AND4 (N9444, N9442, N4001, N9432, N5060);
nor NOR4 (N9445, N2260, N6152, N8391, N2390);
and AND4 (N9446, N9437, N1995, N1366, N7569);
buf BUF1 (N9447, N9445);
xor XOR2 (N9448, N9447, N8117);
nand NAND4 (N9449, N9446, N1360, N884, N7612);
or OR2 (N9450, N9440, N203);
or OR3 (N9451, N9441, N1131, N5467);
nor NOR2 (N9452, N9431, N2349);
or OR2 (N9453, N9438, N9272);
nor NOR2 (N9454, N9452, N3851);
nand NAND4 (N9455, N9443, N9202, N4803, N1438);
not NOT1 (N9456, N9451);
nand NAND4 (N9457, N9453, N2912, N3085, N2632);
nor NOR4 (N9458, N9444, N4064, N5983, N657);
and AND2 (N9459, N9434, N4281);
nor NOR2 (N9460, N9459, N3428);
not NOT1 (N9461, N9450);
xor XOR2 (N9462, N9461, N4093);
or OR3 (N9463, N9449, N2963, N379);
xor XOR2 (N9464, N9457, N5612);
not NOT1 (N9465, N9458);
nand NAND3 (N9466, N9460, N7068, N309);
nand NAND4 (N9467, N9466, N6383, N7399, N1598);
nor NOR2 (N9468, N9467, N4606);
nand NAND4 (N9469, N9455, N7441, N9397, N136);
nor NOR2 (N9470, N9469, N4165);
buf BUF1 (N9471, N9463);
xor XOR2 (N9472, N9454, N1534);
or OR2 (N9473, N9468, N5820);
nor NOR4 (N9474, N9471, N6911, N3446, N3061);
nand NAND3 (N9475, N9474, N9314, N7812);
xor XOR2 (N9476, N9470, N1846);
nand NAND2 (N9477, N9448, N6159);
or OR4 (N9478, N9475, N6853, N2102, N1120);
not NOT1 (N9479, N9473);
xor XOR2 (N9480, N9476, N7410);
xor XOR2 (N9481, N9477, N3742);
buf BUF1 (N9482, N9464);
and AND3 (N9483, N9480, N4429, N2631);
and AND3 (N9484, N9479, N1266, N5230);
nand NAND3 (N9485, N9482, N3512, N8918);
not NOT1 (N9486, N9456);
or OR2 (N9487, N9435, N6413);
and AND4 (N9488, N9483, N5823, N9482, N2202);
or OR4 (N9489, N9486, N2733, N9225, N6539);
and AND3 (N9490, N9481, N9448, N2792);
not NOT1 (N9491, N9484);
or OR4 (N9492, N9490, N4326, N6738, N2823);
nand NAND3 (N9493, N9472, N7222, N1662);
buf BUF1 (N9494, N9465);
buf BUF1 (N9495, N9485);
not NOT1 (N9496, N9495);
and AND2 (N9497, N9494, N413);
nor NOR3 (N9498, N9493, N1992, N6709);
nand NAND3 (N9499, N9498, N1342, N9461);
nand NAND4 (N9500, N9491, N2367, N3643, N3926);
xor XOR2 (N9501, N9489, N7371);
not NOT1 (N9502, N9497);
nor NOR2 (N9503, N9492, N3230);
or OR4 (N9504, N9462, N6733, N6572, N9210);
and AND4 (N9505, N9501, N1275, N3199, N3499);
buf BUF1 (N9506, N9503);
not NOT1 (N9507, N9488);
or OR3 (N9508, N9502, N9088, N7651);
or OR3 (N9509, N9504, N7793, N2770);
and AND3 (N9510, N9496, N6561, N9444);
not NOT1 (N9511, N9508);
and AND3 (N9512, N9505, N3965, N4679);
or OR4 (N9513, N9507, N1088, N2316, N8228);
not NOT1 (N9514, N9478);
or OR3 (N9515, N9513, N7112, N4828);
and AND4 (N9516, N9506, N5921, N2768, N4853);
and AND3 (N9517, N9514, N2758, N9423);
not NOT1 (N9518, N9515);
and AND3 (N9519, N9499, N1211, N8630);
or OR4 (N9520, N9487, N917, N5983, N9266);
buf BUF1 (N9521, N9518);
not NOT1 (N9522, N9511);
nand NAND4 (N9523, N9512, N6722, N3947, N1076);
buf BUF1 (N9524, N9521);
and AND2 (N9525, N9524, N2576);
buf BUF1 (N9526, N9509);
and AND2 (N9527, N9523, N2397);
nand NAND4 (N9528, N9517, N9005, N1971, N4218);
and AND4 (N9529, N9528, N1252, N7658, N3543);
buf BUF1 (N9530, N9527);
nor NOR3 (N9531, N9529, N8001, N7523);
buf BUF1 (N9532, N9522);
buf BUF1 (N9533, N9520);
and AND2 (N9534, N9531, N4511);
buf BUF1 (N9535, N9500);
not NOT1 (N9536, N9533);
xor XOR2 (N9537, N9510, N5645);
not NOT1 (N9538, N9535);
not NOT1 (N9539, N9536);
not NOT1 (N9540, N9532);
buf BUF1 (N9541, N9525);
not NOT1 (N9542, N9519);
nor NOR4 (N9543, N9541, N1551, N3927, N6806);
and AND2 (N9544, N9539, N3876);
buf BUF1 (N9545, N9542);
nand NAND2 (N9546, N9516, N116);
nand NAND3 (N9547, N9534, N1835, N2771);
buf BUF1 (N9548, N9530);
not NOT1 (N9549, N9544);
or OR2 (N9550, N9547, N887);
xor XOR2 (N9551, N9546, N5166);
or OR3 (N9552, N9543, N1534, N5879);
or OR3 (N9553, N9550, N3943, N8448);
xor XOR2 (N9554, N9540, N6285);
nand NAND4 (N9555, N9554, N3174, N4397, N632);
nor NOR4 (N9556, N9526, N8006, N1406, N3792);
nand NAND3 (N9557, N9552, N2418, N7804);
xor XOR2 (N9558, N9548, N1855);
nor NOR4 (N9559, N9555, N5671, N2721, N4986);
buf BUF1 (N9560, N9556);
or OR4 (N9561, N9545, N7462, N1715, N4291);
nand NAND3 (N9562, N9559, N861, N5778);
xor XOR2 (N9563, N9551, N2941);
xor XOR2 (N9564, N9561, N3658);
nor NOR3 (N9565, N9560, N6610, N1105);
nor NOR4 (N9566, N9553, N1513, N2960, N2414);
not NOT1 (N9567, N9565);
nand NAND3 (N9568, N9537, N6447, N7864);
buf BUF1 (N9569, N9558);
and AND3 (N9570, N9549, N8932, N7524);
and AND3 (N9571, N9570, N6959, N6806);
nor NOR2 (N9572, N9538, N3179);
xor XOR2 (N9573, N9562, N3857);
or OR4 (N9574, N9567, N1438, N3377, N4573);
buf BUF1 (N9575, N9568);
or OR4 (N9576, N9563, N8024, N7588, N2306);
nand NAND3 (N9577, N9574, N248, N8725);
or OR4 (N9578, N9577, N8199, N6942, N8907);
nor NOR3 (N9579, N9575, N6103, N9077);
or OR3 (N9580, N9571, N6589, N9238);
not NOT1 (N9581, N9572);
nor NOR4 (N9582, N9557, N3003, N9405, N7730);
xor XOR2 (N9583, N9564, N3896);
buf BUF1 (N9584, N9566);
or OR2 (N9585, N9580, N1961);
nor NOR2 (N9586, N9581, N773);
buf BUF1 (N9587, N9579);
and AND4 (N9588, N9586, N1377, N5175, N5105);
or OR3 (N9589, N9573, N4779, N3899);
and AND3 (N9590, N9584, N4444, N2418);
and AND3 (N9591, N9589, N7855, N5783);
nand NAND4 (N9592, N9591, N8965, N2456, N7052);
xor XOR2 (N9593, N9583, N5342);
or OR4 (N9594, N9588, N7985, N1417, N1077);
not NOT1 (N9595, N9569);
buf BUF1 (N9596, N9590);
nor NOR3 (N9597, N9592, N1472, N6958);
not NOT1 (N9598, N9587);
xor XOR2 (N9599, N9576, N1121);
buf BUF1 (N9600, N9594);
and AND2 (N9601, N9582, N7470);
buf BUF1 (N9602, N9585);
nand NAND4 (N9603, N9595, N5456, N7381, N657);
nand NAND2 (N9604, N9597, N7766);
not NOT1 (N9605, N9596);
xor XOR2 (N9606, N9593, N2030);
and AND4 (N9607, N9602, N6568, N828, N3101);
xor XOR2 (N9608, N9603, N482);
or OR3 (N9609, N9607, N8562, N4628);
not NOT1 (N9610, N9599);
xor XOR2 (N9611, N9601, N6302);
xor XOR2 (N9612, N9605, N3300);
nand NAND2 (N9613, N9606, N2236);
nand NAND3 (N9614, N9598, N8020, N1434);
and AND3 (N9615, N9612, N6271, N9505);
not NOT1 (N9616, N9604);
and AND2 (N9617, N9610, N8339);
not NOT1 (N9618, N9600);
nand NAND4 (N9619, N9614, N7160, N3079, N5679);
xor XOR2 (N9620, N9619, N6107);
xor XOR2 (N9621, N9618, N6148);
nor NOR4 (N9622, N9578, N8103, N7315, N3329);
nand NAND3 (N9623, N9617, N1386, N8565);
buf BUF1 (N9624, N9608);
xor XOR2 (N9625, N9611, N9574);
nand NAND2 (N9626, N9613, N5694);
and AND3 (N9627, N9626, N1893, N2616);
and AND3 (N9628, N9623, N6100, N1745);
not NOT1 (N9629, N9628);
xor XOR2 (N9630, N9609, N9052);
nor NOR2 (N9631, N9629, N5662);
and AND4 (N9632, N9621, N742, N9163, N5337);
xor XOR2 (N9633, N9620, N1252);
nand NAND4 (N9634, N9632, N5338, N7006, N7566);
buf BUF1 (N9635, N9634);
and AND3 (N9636, N9616, N8006, N5173);
or OR2 (N9637, N9630, N8616);
or OR3 (N9638, N9631, N3409, N4443);
nor NOR3 (N9639, N9638, N5898, N2110);
nand NAND2 (N9640, N9639, N707);
buf BUF1 (N9641, N9622);
not NOT1 (N9642, N9641);
buf BUF1 (N9643, N9625);
nand NAND4 (N9644, N9637, N9514, N4603, N9138);
buf BUF1 (N9645, N9636);
and AND4 (N9646, N9633, N8389, N2222, N7401);
and AND3 (N9647, N9624, N3085, N2138);
or OR4 (N9648, N9615, N2192, N8023, N204);
buf BUF1 (N9649, N9644);
xor XOR2 (N9650, N9646, N6535);
nor NOR4 (N9651, N9650, N4267, N1436, N5835);
nand NAND3 (N9652, N9647, N9063, N1336);
and AND4 (N9653, N9640, N7659, N1037, N7405);
xor XOR2 (N9654, N9649, N4546);
not NOT1 (N9655, N9635);
or OR2 (N9656, N9655, N1345);
buf BUF1 (N9657, N9642);
and AND4 (N9658, N9627, N1922, N922, N7951);
buf BUF1 (N9659, N9651);
not NOT1 (N9660, N9653);
buf BUF1 (N9661, N9658);
buf BUF1 (N9662, N9643);
and AND2 (N9663, N9660, N2780);
xor XOR2 (N9664, N9659, N2075);
or OR2 (N9665, N9662, N2749);
and AND3 (N9666, N9657, N3396, N522);
nand NAND2 (N9667, N9665, N5423);
xor XOR2 (N9668, N9663, N7791);
nand NAND2 (N9669, N9654, N7373);
not NOT1 (N9670, N9667);
not NOT1 (N9671, N9656);
or OR3 (N9672, N9664, N382, N5760);
nand NAND3 (N9673, N9669, N4701, N3083);
or OR4 (N9674, N9673, N3113, N1324, N1248);
and AND2 (N9675, N9668, N6656);
not NOT1 (N9676, N9674);
xor XOR2 (N9677, N9672, N1376);
nor NOR2 (N9678, N9652, N2516);
nand NAND3 (N9679, N9661, N3202, N9513);
and AND3 (N9680, N9671, N2144, N1931);
buf BUF1 (N9681, N9680);
buf BUF1 (N9682, N9666);
nor NOR4 (N9683, N9681, N4771, N2454, N3227);
nand NAND4 (N9684, N9683, N2742, N3825, N1016);
not NOT1 (N9685, N9675);
nand NAND4 (N9686, N9679, N2115, N2780, N8940);
nand NAND2 (N9687, N9684, N7596);
nand NAND2 (N9688, N9685, N4467);
and AND2 (N9689, N9677, N6072);
nand NAND2 (N9690, N9682, N1309);
and AND2 (N9691, N9690, N1200);
or OR4 (N9692, N9689, N1405, N5540, N9670);
or OR3 (N9693, N3627, N3479, N4920);
xor XOR2 (N9694, N9692, N2569);
or OR3 (N9695, N9693, N4165, N7362);
or OR2 (N9696, N9695, N4229);
buf BUF1 (N9697, N9696);
or OR3 (N9698, N9676, N7055, N1635);
or OR4 (N9699, N9691, N8120, N3674, N6728);
or OR3 (N9700, N9694, N7802, N2163);
xor XOR2 (N9701, N9688, N8295);
and AND2 (N9702, N9700, N8192);
and AND2 (N9703, N9678, N6368);
or OR4 (N9704, N9687, N1076, N5582, N3461);
nor NOR3 (N9705, N9704, N2404, N5238);
buf BUF1 (N9706, N9705);
xor XOR2 (N9707, N9686, N7131);
buf BUF1 (N9708, N9645);
not NOT1 (N9709, N9702);
nand NAND3 (N9710, N9697, N864, N358);
nor NOR3 (N9711, N9707, N818, N7518);
nor NOR2 (N9712, N9709, N2685);
and AND3 (N9713, N9710, N7739, N7165);
xor XOR2 (N9714, N9706, N642);
nor NOR2 (N9715, N9699, N4975);
buf BUF1 (N9716, N9715);
and AND3 (N9717, N9716, N5662, N9131);
nand NAND4 (N9718, N9717, N3889, N4289, N6770);
nor NOR3 (N9719, N9698, N694, N7797);
nor NOR2 (N9720, N9719, N3865);
nor NOR4 (N9721, N9713, N8152, N5352, N2392);
nand NAND3 (N9722, N9718, N3466, N2400);
or OR4 (N9723, N9711, N6274, N2901, N2565);
not NOT1 (N9724, N9648);
and AND4 (N9725, N9703, N1587, N4393, N4719);
or OR2 (N9726, N9721, N8686);
or OR2 (N9727, N9725, N746);
and AND2 (N9728, N9708, N2871);
not NOT1 (N9729, N9727);
not NOT1 (N9730, N9722);
nand NAND2 (N9731, N9701, N706);
xor XOR2 (N9732, N9714, N3074);
xor XOR2 (N9733, N9724, N1219);
buf BUF1 (N9734, N9730);
xor XOR2 (N9735, N9732, N1867);
nand NAND4 (N9736, N9733, N4006, N6080, N2051);
buf BUF1 (N9737, N9734);
nand NAND2 (N9738, N9723, N7227);
buf BUF1 (N9739, N9738);
nor NOR3 (N9740, N9737, N1210, N4805);
nand NAND4 (N9741, N9720, N1617, N6144, N5916);
and AND2 (N9742, N9741, N1635);
nor NOR4 (N9743, N9740, N6559, N8147, N9499);
and AND3 (N9744, N9739, N7539, N7418);
or OR4 (N9745, N9742, N709, N7119, N3690);
buf BUF1 (N9746, N9744);
not NOT1 (N9747, N9735);
nor NOR4 (N9748, N9712, N8319, N6666, N6479);
xor XOR2 (N9749, N9743, N461);
xor XOR2 (N9750, N9746, N3134);
buf BUF1 (N9751, N9731);
or OR2 (N9752, N9749, N7180);
and AND4 (N9753, N9748, N3017, N3368, N5392);
or OR3 (N9754, N9752, N8051, N5435);
xor XOR2 (N9755, N9751, N4825);
not NOT1 (N9756, N9750);
xor XOR2 (N9757, N9755, N3253);
or OR4 (N9758, N9756, N7196, N8175, N3775);
or OR2 (N9759, N9729, N5182);
nor NOR3 (N9760, N9726, N7769, N6574);
xor XOR2 (N9761, N9759, N1430);
buf BUF1 (N9762, N9761);
nor NOR4 (N9763, N9757, N4826, N3880, N3226);
and AND4 (N9764, N9747, N8294, N6176, N3876);
xor XOR2 (N9765, N9745, N465);
nand NAND3 (N9766, N9758, N7345, N5898);
not NOT1 (N9767, N9766);
nand NAND4 (N9768, N9760, N4526, N1898, N4974);
xor XOR2 (N9769, N9736, N565);
nor NOR4 (N9770, N9767, N7718, N5546, N6098);
buf BUF1 (N9771, N9768);
or OR4 (N9772, N9769, N4809, N9160, N1916);
nand NAND3 (N9773, N9765, N4853, N7758);
nor NOR2 (N9774, N9762, N2654);
buf BUF1 (N9775, N9771);
buf BUF1 (N9776, N9728);
and AND3 (N9777, N9770, N5028, N6909);
xor XOR2 (N9778, N9775, N9435);
xor XOR2 (N9779, N9774, N7722);
not NOT1 (N9780, N9764);
not NOT1 (N9781, N9772);
nor NOR4 (N9782, N9773, N4001, N8865, N3131);
or OR3 (N9783, N9753, N8980, N7437);
nor NOR3 (N9784, N9780, N8883, N8675);
nor NOR3 (N9785, N9763, N4558, N1300);
xor XOR2 (N9786, N9754, N8960);
nand NAND4 (N9787, N9782, N9141, N4782, N3273);
xor XOR2 (N9788, N9779, N8733);
and AND4 (N9789, N9787, N1627, N2052, N1997);
and AND3 (N9790, N9777, N105, N1398);
xor XOR2 (N9791, N9784, N3801);
not NOT1 (N9792, N9790);
and AND3 (N9793, N9778, N9748, N5119);
nor NOR4 (N9794, N9792, N6762, N5378, N9765);
not NOT1 (N9795, N9786);
or OR2 (N9796, N9789, N7341);
nand NAND4 (N9797, N9796, N6403, N6465, N185);
xor XOR2 (N9798, N9788, N838);
nand NAND3 (N9799, N9783, N4928, N3588);
nor NOR4 (N9800, N9776, N576, N5641, N1195);
not NOT1 (N9801, N9798);
buf BUF1 (N9802, N9797);
or OR2 (N9803, N9802, N9161);
or OR3 (N9804, N9785, N4421, N6486);
not NOT1 (N9805, N9781);
buf BUF1 (N9806, N9803);
nor NOR3 (N9807, N9801, N7008, N8264);
buf BUF1 (N9808, N9791);
xor XOR2 (N9809, N9805, N184);
or OR4 (N9810, N9793, N706, N4436, N364);
xor XOR2 (N9811, N9806, N9588);
xor XOR2 (N9812, N9811, N478);
xor XOR2 (N9813, N9800, N6592);
not NOT1 (N9814, N9794);
not NOT1 (N9815, N9812);
nor NOR4 (N9816, N9813, N1083, N5975, N8176);
not NOT1 (N9817, N9815);
xor XOR2 (N9818, N9799, N8862);
buf BUF1 (N9819, N9807);
and AND3 (N9820, N9818, N1137, N2241);
nor NOR4 (N9821, N9810, N1798, N8921, N3004);
nand NAND3 (N9822, N9809, N4783, N8081);
not NOT1 (N9823, N9821);
or OR4 (N9824, N9816, N1588, N7079, N7142);
or OR3 (N9825, N9822, N3355, N4573);
xor XOR2 (N9826, N9804, N8332);
or OR3 (N9827, N9817, N9420, N5539);
nor NOR4 (N9828, N9795, N1535, N9608, N6079);
not NOT1 (N9829, N9826);
and AND2 (N9830, N9825, N944);
xor XOR2 (N9831, N9828, N9366);
or OR2 (N9832, N9829, N2092);
nor NOR2 (N9833, N9823, N8859);
or OR2 (N9834, N9831, N3193);
or OR2 (N9835, N9827, N8573);
buf BUF1 (N9836, N9824);
or OR3 (N9837, N9808, N3651, N8981);
xor XOR2 (N9838, N9834, N5392);
nor NOR3 (N9839, N9836, N1858, N2336);
xor XOR2 (N9840, N9820, N8217);
or OR2 (N9841, N9838, N9208);
nand NAND4 (N9842, N9830, N6873, N4789, N4460);
nor NOR2 (N9843, N9840, N4057);
nand NAND4 (N9844, N9819, N4722, N706, N2228);
and AND3 (N9845, N9839, N3180, N2899);
not NOT1 (N9846, N9842);
buf BUF1 (N9847, N9844);
xor XOR2 (N9848, N9845, N3538);
xor XOR2 (N9849, N9848, N5324);
buf BUF1 (N9850, N9832);
or OR3 (N9851, N9837, N9776, N1446);
xor XOR2 (N9852, N9849, N1127);
buf BUF1 (N9853, N9843);
and AND3 (N9854, N9853, N9740, N2262);
xor XOR2 (N9855, N9851, N5698);
nor NOR2 (N9856, N9852, N7904);
nand NAND3 (N9857, N9854, N5795, N1058);
and AND3 (N9858, N9847, N8272, N4157);
and AND2 (N9859, N9855, N2469);
nor NOR3 (N9860, N9858, N8127, N5266);
not NOT1 (N9861, N9859);
nor NOR2 (N9862, N9846, N4094);
xor XOR2 (N9863, N9814, N3979);
nand NAND2 (N9864, N9850, N9190);
nor NOR3 (N9865, N9860, N3178, N1104);
buf BUF1 (N9866, N9864);
or OR2 (N9867, N9863, N5872);
nand NAND4 (N9868, N9861, N1384, N8919, N3014);
or OR2 (N9869, N9835, N3635);
not NOT1 (N9870, N9841);
and AND4 (N9871, N9862, N3152, N3583, N994);
and AND4 (N9872, N9866, N1387, N7683, N3282);
not NOT1 (N9873, N9868);
not NOT1 (N9874, N9833);
xor XOR2 (N9875, N9856, N8398);
xor XOR2 (N9876, N9874, N8337);
nor NOR4 (N9877, N9873, N2630, N5505, N9653);
nand NAND4 (N9878, N9877, N9114, N9422, N3930);
xor XOR2 (N9879, N9857, N573);
not NOT1 (N9880, N9865);
not NOT1 (N9881, N9876);
not NOT1 (N9882, N9881);
nand NAND4 (N9883, N9869, N7209, N115, N7127);
not NOT1 (N9884, N9879);
not NOT1 (N9885, N9870);
or OR2 (N9886, N9885, N2429);
nor NOR2 (N9887, N9886, N4642);
nand NAND4 (N9888, N9872, N8456, N8975, N1521);
buf BUF1 (N9889, N9867);
nor NOR4 (N9890, N9882, N7954, N3208, N2256);
or OR3 (N9891, N9884, N5939, N8819);
or OR4 (N9892, N9888, N2490, N8255, N6578);
nand NAND2 (N9893, N9887, N9676);
not NOT1 (N9894, N9890);
not NOT1 (N9895, N9883);
and AND4 (N9896, N9895, N6569, N2536, N6101);
buf BUF1 (N9897, N9889);
not NOT1 (N9898, N9880);
not NOT1 (N9899, N9878);
or OR2 (N9900, N9875, N3010);
and AND3 (N9901, N9898, N7906, N4792);
buf BUF1 (N9902, N9897);
nor NOR4 (N9903, N9894, N4537, N823, N1585);
buf BUF1 (N9904, N9902);
nand NAND4 (N9905, N9871, N4127, N2803, N4691);
xor XOR2 (N9906, N9904, N5240);
nand NAND2 (N9907, N9900, N3905);
or OR2 (N9908, N9899, N1486);
not NOT1 (N9909, N9905);
nor NOR2 (N9910, N9901, N2267);
nor NOR2 (N9911, N9908, N541);
buf BUF1 (N9912, N9907);
xor XOR2 (N9913, N9906, N3495);
xor XOR2 (N9914, N9893, N7894);
nand NAND2 (N9915, N9913, N5871);
xor XOR2 (N9916, N9911, N9428);
or OR4 (N9917, N9912, N5883, N2866, N5534);
nand NAND3 (N9918, N9903, N7076, N6137);
xor XOR2 (N9919, N9915, N6471);
xor XOR2 (N9920, N9918, N199);
buf BUF1 (N9921, N9917);
and AND2 (N9922, N9914, N8309);
nor NOR4 (N9923, N9919, N3106, N9390, N5685);
nand NAND4 (N9924, N9891, N9904, N2535, N8024);
buf BUF1 (N9925, N9924);
nor NOR4 (N9926, N9896, N457, N9486, N7411);
not NOT1 (N9927, N9925);
not NOT1 (N9928, N9920);
not NOT1 (N9929, N9922);
buf BUF1 (N9930, N9926);
nand NAND4 (N9931, N9927, N6201, N746, N5276);
not NOT1 (N9932, N9916);
buf BUF1 (N9933, N9909);
or OR3 (N9934, N9932, N1750, N9651);
xor XOR2 (N9935, N9931, N7249);
or OR2 (N9936, N9930, N3934);
xor XOR2 (N9937, N9892, N775);
and AND2 (N9938, N9937, N7879);
not NOT1 (N9939, N9935);
or OR4 (N9940, N9936, N9683, N9478, N666);
xor XOR2 (N9941, N9933, N897);
not NOT1 (N9942, N9939);
buf BUF1 (N9943, N9921);
or OR3 (N9944, N9928, N3270, N9758);
nor NOR3 (N9945, N9929, N4518, N113);
nor NOR4 (N9946, N9910, N5823, N1309, N199);
nand NAND4 (N9947, N9941, N1373, N3901, N3251);
not NOT1 (N9948, N9945);
or OR3 (N9949, N9948, N3618, N5419);
nand NAND4 (N9950, N9934, N9783, N537, N5870);
nand NAND2 (N9951, N9946, N5270);
nor NOR3 (N9952, N9938, N7042, N3302);
nand NAND3 (N9953, N9943, N7423, N5352);
nor NOR2 (N9954, N9952, N4655);
or OR2 (N9955, N9953, N2915);
xor XOR2 (N9956, N9949, N3949);
xor XOR2 (N9957, N9942, N2270);
and AND4 (N9958, N9950, N2704, N5499, N6683);
xor XOR2 (N9959, N9954, N2668);
and AND3 (N9960, N9958, N3356, N4096);
nand NAND4 (N9961, N9955, N2837, N8825, N2452);
or OR3 (N9962, N9944, N5563, N7518);
not NOT1 (N9963, N9960);
or OR2 (N9964, N9940, N5837);
and AND4 (N9965, N9964, N1420, N9888, N2647);
buf BUF1 (N9966, N9961);
buf BUF1 (N9967, N9963);
nor NOR3 (N9968, N9951, N8024, N3537);
not NOT1 (N9969, N9965);
or OR4 (N9970, N9959, N7299, N2398, N4510);
and AND3 (N9971, N9969, N5475, N8163);
not NOT1 (N9972, N9923);
or OR4 (N9973, N9970, N919, N6926, N9424);
or OR4 (N9974, N9962, N8591, N3661, N3311);
nand NAND4 (N9975, N9973, N5976, N649, N3898);
not NOT1 (N9976, N9971);
nand NAND2 (N9977, N9974, N5061);
xor XOR2 (N9978, N9966, N2586);
buf BUF1 (N9979, N9972);
nor NOR2 (N9980, N9979, N381);
and AND4 (N9981, N9957, N3016, N1654, N4552);
not NOT1 (N9982, N9968);
not NOT1 (N9983, N9980);
and AND4 (N9984, N9947, N2814, N3474, N5199);
or OR3 (N9985, N9967, N7167, N4062);
buf BUF1 (N9986, N9983);
nor NOR3 (N9987, N9956, N2684, N8233);
nor NOR4 (N9988, N9986, N5585, N1139, N4264);
and AND2 (N9989, N9978, N9237);
nor NOR4 (N9990, N9987, N8881, N4405, N3234);
not NOT1 (N9991, N9975);
or OR2 (N9992, N9990, N2925);
xor XOR2 (N9993, N9977, N3603);
xor XOR2 (N9994, N9991, N7918);
not NOT1 (N9995, N9982);
or OR3 (N9996, N9985, N5646, N8119);
nand NAND2 (N9997, N9988, N7023);
nor NOR4 (N9998, N9995, N5138, N2054, N1167);
and AND3 (N9999, N9989, N2109, N3108);
and AND2 (N10000, N9976, N2374);
or OR2 (N10001, N9994, N7679);
not NOT1 (N10002, N9981);
xor XOR2 (N10003, N9984, N8417);
buf BUF1 (N10004, N10002);
nor NOR3 (N10005, N9998, N5966, N6165);
nor NOR3 (N10006, N10000, N4335, N8784);
xor XOR2 (N10007, N10006, N8557);
not NOT1 (N10008, N10003);
nor NOR2 (N10009, N9993, N1749);
or OR2 (N10010, N10009, N6487);
and AND2 (N10011, N9996, N2241);
buf BUF1 (N10012, N10008);
not NOT1 (N10013, N10001);
or OR3 (N10014, N9999, N7238, N8935);
or OR2 (N10015, N10014, N4079);
nor NOR4 (N10016, N10007, N9581, N4793, N979);
and AND3 (N10017, N10016, N2856, N9417);
nor NOR2 (N10018, N10013, N2316);
nand NAND4 (N10019, N9997, N6247, N7804, N5106);
xor XOR2 (N10020, N10019, N8908);
not NOT1 (N10021, N10012);
nand NAND2 (N10022, N10004, N7779);
buf BUF1 (N10023, N10017);
nand NAND4 (N10024, N10005, N4623, N1268, N26);
and AND4 (N10025, N10024, N7862, N9795, N6850);
nor NOR3 (N10026, N10015, N1568, N6927);
not NOT1 (N10027, N9992);
and AND4 (N10028, N10010, N2332, N6237, N2044);
or OR2 (N10029, N10025, N6715);
nand NAND4 (N10030, N10020, N5768, N6990, N8677);
nor NOR2 (N10031, N10028, N8089);
and AND2 (N10032, N10021, N3672);
buf BUF1 (N10033, N10018);
buf BUF1 (N10034, N10030);
and AND3 (N10035, N10033, N7259, N3136);
buf BUF1 (N10036, N10023);
not NOT1 (N10037, N10011);
and AND4 (N10038, N10037, N9869, N4142, N2203);
not NOT1 (N10039, N10026);
not NOT1 (N10040, N10036);
nand NAND4 (N10041, N10031, N3938, N8051, N5438);
or OR2 (N10042, N10035, N7497);
or OR4 (N10043, N10032, N2116, N4658, N8269);
xor XOR2 (N10044, N10041, N6666);
and AND3 (N10045, N10029, N3130, N5211);
nand NAND3 (N10046, N10039, N8247, N2337);
and AND4 (N10047, N10038, N6394, N3076, N2227);
nor NOR3 (N10048, N10044, N6408, N3923);
nand NAND3 (N10049, N10022, N6379, N4615);
nand NAND2 (N10050, N10040, N512);
not NOT1 (N10051, N10043);
nand NAND4 (N10052, N10034, N7110, N475, N7836);
nor NOR4 (N10053, N10051, N9570, N9427, N3068);
nor NOR2 (N10054, N10048, N2584);
nor NOR2 (N10055, N10047, N7412);
not NOT1 (N10056, N10046);
buf BUF1 (N10057, N10053);
xor XOR2 (N10058, N10050, N9155);
xor XOR2 (N10059, N10055, N5116);
nand NAND2 (N10060, N10057, N7901);
not NOT1 (N10061, N10056);
or OR3 (N10062, N10042, N3860, N3059);
nor NOR4 (N10063, N10054, N3917, N8230, N4690);
not NOT1 (N10064, N10027);
nor NOR4 (N10065, N10059, N3083, N3700, N2641);
not NOT1 (N10066, N10065);
not NOT1 (N10067, N10062);
nand NAND2 (N10068, N10067, N9720);
nand NAND4 (N10069, N10063, N9603, N1766, N4942);
not NOT1 (N10070, N10064);
or OR4 (N10071, N10066, N5592, N4262, N5745);
or OR2 (N10072, N10049, N8841);
or OR4 (N10073, N10071, N9176, N4986, N2567);
xor XOR2 (N10074, N10073, N2736);
nor NOR2 (N10075, N10060, N1375);
and AND2 (N10076, N10061, N2374);
or OR2 (N10077, N10072, N5219);
or OR4 (N10078, N10070, N6706, N8950, N2124);
or OR2 (N10079, N10076, N2416);
buf BUF1 (N10080, N10068);
or OR2 (N10081, N10078, N8413);
nor NOR4 (N10082, N10075, N1988, N7512, N8916);
nor NOR3 (N10083, N10077, N7297, N3552);
xor XOR2 (N10084, N10058, N4171);
or OR4 (N10085, N10083, N2344, N877, N2483);
and AND3 (N10086, N10085, N8233, N9684);
nand NAND3 (N10087, N10069, N5466, N8970);
buf BUF1 (N10088, N10079);
and AND4 (N10089, N10074, N6085, N5897, N7943);
and AND4 (N10090, N10045, N4778, N8782, N926);
nor NOR4 (N10091, N10089, N3354, N10065, N1075);
or OR4 (N10092, N10082, N9929, N31, N3425);
buf BUF1 (N10093, N10080);
nand NAND2 (N10094, N10086, N9547);
nand NAND3 (N10095, N10081, N368, N7884);
nand NAND3 (N10096, N10094, N874, N404);
buf BUF1 (N10097, N10091);
xor XOR2 (N10098, N10095, N6274);
nor NOR4 (N10099, N10092, N185, N1174, N2208);
nand NAND4 (N10100, N10087, N6388, N4777, N2963);
and AND3 (N10101, N10090, N8082, N7014);
xor XOR2 (N10102, N10084, N7443);
and AND3 (N10103, N10097, N7355, N3167);
or OR3 (N10104, N10100, N4901, N5272);
buf BUF1 (N10105, N10099);
nor NOR4 (N10106, N10093, N9914, N5037, N4666);
nor NOR4 (N10107, N10102, N3818, N10093, N5443);
nor NOR3 (N10108, N10096, N2953, N387);
buf BUF1 (N10109, N10107);
nand NAND2 (N10110, N10105, N4611);
buf BUF1 (N10111, N10109);
or OR2 (N10112, N10106, N2208);
buf BUF1 (N10113, N10101);
nor NOR2 (N10114, N10111, N3680);
not NOT1 (N10115, N10112);
nor NOR4 (N10116, N10114, N5861, N8449, N9651);
xor XOR2 (N10117, N10104, N3269);
xor XOR2 (N10118, N10098, N3875);
buf BUF1 (N10119, N10088);
and AND4 (N10120, N10113, N2701, N4144, N7172);
buf BUF1 (N10121, N10103);
and AND3 (N10122, N10052, N1069, N6809);
not NOT1 (N10123, N10121);
nor NOR3 (N10124, N10108, N6004, N6131);
buf BUF1 (N10125, N10119);
and AND2 (N10126, N10115, N3833);
buf BUF1 (N10127, N10124);
and AND4 (N10128, N10110, N2580, N920, N5789);
not NOT1 (N10129, N10127);
xor XOR2 (N10130, N10116, N6466);
xor XOR2 (N10131, N10125, N4274);
nor NOR4 (N10132, N10123, N5482, N2657, N5318);
or OR2 (N10133, N10130, N1660);
xor XOR2 (N10134, N10131, N5265);
and AND3 (N10135, N10122, N111, N5677);
nor NOR4 (N10136, N10134, N8811, N4475, N6758);
and AND2 (N10137, N10117, N503);
buf BUF1 (N10138, N10126);
not NOT1 (N10139, N10129);
xor XOR2 (N10140, N10135, N6324);
nor NOR3 (N10141, N10118, N1999, N4439);
nor NOR3 (N10142, N10141, N6708, N627);
xor XOR2 (N10143, N10132, N895);
not NOT1 (N10144, N10139);
or OR3 (N10145, N10140, N9920, N2631);
buf BUF1 (N10146, N10142);
nor NOR2 (N10147, N10133, N4791);
not NOT1 (N10148, N10138);
and AND3 (N10149, N10145, N6257, N4925);
not NOT1 (N10150, N10148);
nand NAND4 (N10151, N10137, N7758, N3418, N9502);
not NOT1 (N10152, N10143);
or OR4 (N10153, N10150, N7124, N8221, N9736);
nand NAND4 (N10154, N10149, N5865, N5555, N7802);
not NOT1 (N10155, N10147);
buf BUF1 (N10156, N10153);
buf BUF1 (N10157, N10120);
xor XOR2 (N10158, N10151, N5392);
and AND4 (N10159, N10144, N4403, N1731, N9936);
not NOT1 (N10160, N10136);
and AND2 (N10161, N10157, N7011);
or OR3 (N10162, N10161, N8938, N3063);
or OR2 (N10163, N10160, N5033);
buf BUF1 (N10164, N10128);
or OR3 (N10165, N10159, N7998, N4453);
or OR3 (N10166, N10156, N9166, N8563);
xor XOR2 (N10167, N10154, N1765);
xor XOR2 (N10168, N10164, N8812);
xor XOR2 (N10169, N10165, N2244);
buf BUF1 (N10170, N10152);
or OR2 (N10171, N10162, N1122);
buf BUF1 (N10172, N10158);
and AND2 (N10173, N10146, N8607);
nor NOR3 (N10174, N10171, N7435, N700);
and AND4 (N10175, N10169, N3838, N8025, N9977);
buf BUF1 (N10176, N10173);
or OR2 (N10177, N10170, N6351);
nand NAND2 (N10178, N10168, N7092);
xor XOR2 (N10179, N10163, N6513);
or OR3 (N10180, N10172, N1411, N8406);
not NOT1 (N10181, N10155);
nor NOR2 (N10182, N10178, N6577);
xor XOR2 (N10183, N10180, N478);
not NOT1 (N10184, N10174);
nand NAND3 (N10185, N10182, N8211, N5560);
xor XOR2 (N10186, N10176, N2609);
nand NAND2 (N10187, N10186, N2337);
nor NOR2 (N10188, N10175, N3275);
and AND3 (N10189, N10179, N9421, N10175);
not NOT1 (N10190, N10166);
and AND4 (N10191, N10188, N6468, N9532, N7879);
or OR4 (N10192, N10191, N3520, N6195, N5945);
not NOT1 (N10193, N10177);
nand NAND4 (N10194, N10185, N64, N1, N83);
nand NAND4 (N10195, N10190, N8660, N2819, N3529);
nor NOR3 (N10196, N10195, N609, N7807);
and AND4 (N10197, N10187, N658, N7886, N887);
or OR4 (N10198, N10181, N7854, N381, N6787);
and AND3 (N10199, N10192, N7743, N1755);
nand NAND2 (N10200, N10189, N295);
xor XOR2 (N10201, N10183, N1838);
nand NAND2 (N10202, N10200, N8309);
nor NOR3 (N10203, N10194, N6107, N9582);
nor NOR3 (N10204, N10201, N1915, N1281);
nor NOR2 (N10205, N10204, N2948);
or OR2 (N10206, N10196, N4129);
nor NOR3 (N10207, N10205, N2533, N1821);
not NOT1 (N10208, N10206);
or OR4 (N10209, N10199, N3736, N1865, N7427);
buf BUF1 (N10210, N10184);
or OR4 (N10211, N10198, N8958, N2321, N878);
nand NAND2 (N10212, N10203, N2354);
not NOT1 (N10213, N10212);
nor NOR3 (N10214, N10202, N974, N1887);
xor XOR2 (N10215, N10197, N8961);
nand NAND2 (N10216, N10211, N3794);
nand NAND3 (N10217, N10214, N7392, N2976);
not NOT1 (N10218, N10217);
xor XOR2 (N10219, N10215, N6332);
buf BUF1 (N10220, N10167);
or OR2 (N10221, N10209, N7108);
nand NAND2 (N10222, N10210, N7080);
or OR2 (N10223, N10208, N1420);
not NOT1 (N10224, N10218);
and AND2 (N10225, N10207, N5149);
nand NAND3 (N10226, N10193, N463, N1482);
and AND2 (N10227, N10226, N7780);
nor NOR3 (N10228, N10219, N1773, N8526);
buf BUF1 (N10229, N10224);
not NOT1 (N10230, N10225);
xor XOR2 (N10231, N10223, N7412);
nor NOR4 (N10232, N10216, N5648, N1588, N6320);
not NOT1 (N10233, N10229);
and AND2 (N10234, N10221, N6656);
and AND2 (N10235, N10233, N5841);
or OR4 (N10236, N10232, N10224, N164, N1114);
and AND4 (N10237, N10227, N8679, N506, N9219);
not NOT1 (N10238, N10230);
xor XOR2 (N10239, N10231, N5418);
not NOT1 (N10240, N10228);
xor XOR2 (N10241, N10236, N5825);
nand NAND3 (N10242, N10220, N8232, N4487);
nand NAND4 (N10243, N10235, N2587, N3545, N8343);
not NOT1 (N10244, N10241);
buf BUF1 (N10245, N10240);
not NOT1 (N10246, N10244);
xor XOR2 (N10247, N10242, N10061);
or OR4 (N10248, N10237, N9111, N2543, N3547);
or OR2 (N10249, N10246, N2934);
buf BUF1 (N10250, N10239);
and AND3 (N10251, N10250, N9578, N6663);
or OR4 (N10252, N10213, N1350, N5921, N4102);
or OR2 (N10253, N10238, N4646);
or OR2 (N10254, N10222, N6076);
or OR3 (N10255, N10253, N5504, N4504);
or OR3 (N10256, N10245, N7775, N4381);
nand NAND4 (N10257, N10247, N935, N6726, N7735);
xor XOR2 (N10258, N10243, N6002);
nand NAND3 (N10259, N10256, N1800, N5409);
xor XOR2 (N10260, N10254, N4086);
and AND2 (N10261, N10260, N3978);
or OR2 (N10262, N10248, N4126);
nor NOR3 (N10263, N10255, N6334, N5180);
not NOT1 (N10264, N10261);
buf BUF1 (N10265, N10263);
nand NAND2 (N10266, N10262, N7575);
or OR2 (N10267, N10249, N3507);
xor XOR2 (N10268, N10264, N9337);
or OR4 (N10269, N10268, N9780, N212, N4029);
buf BUF1 (N10270, N10266);
buf BUF1 (N10271, N10270);
not NOT1 (N10272, N10265);
not NOT1 (N10273, N10269);
xor XOR2 (N10274, N10251, N6143);
nand NAND2 (N10275, N10258, N7154);
nand NAND4 (N10276, N10252, N3721, N9291, N2859);
xor XOR2 (N10277, N10272, N7421);
nor NOR4 (N10278, N10271, N4061, N7291, N6857);
or OR2 (N10279, N10276, N2752);
xor XOR2 (N10280, N10259, N8927);
or OR3 (N10281, N10267, N3406, N10052);
not NOT1 (N10282, N10277);
or OR4 (N10283, N10273, N4136, N3117, N7501);
buf BUF1 (N10284, N10282);
buf BUF1 (N10285, N10281);
nand NAND4 (N10286, N10285, N4518, N5967, N1001);
xor XOR2 (N10287, N10275, N7035);
buf BUF1 (N10288, N10283);
or OR2 (N10289, N10284, N839);
xor XOR2 (N10290, N10289, N7146);
nand NAND3 (N10291, N10288, N4370, N4093);
nor NOR3 (N10292, N10234, N7920, N7800);
not NOT1 (N10293, N10257);
not NOT1 (N10294, N10292);
nor NOR3 (N10295, N10293, N9062, N2164);
nor NOR4 (N10296, N10291, N333, N1904, N8334);
nor NOR2 (N10297, N10274, N9649);
or OR4 (N10298, N10278, N452, N1542, N6390);
buf BUF1 (N10299, N10296);
nand NAND3 (N10300, N10297, N7748, N6494);
xor XOR2 (N10301, N10290, N249);
xor XOR2 (N10302, N10279, N4539);
not NOT1 (N10303, N10295);
xor XOR2 (N10304, N10301, N2972);
nand NAND2 (N10305, N10304, N6594);
buf BUF1 (N10306, N10302);
not NOT1 (N10307, N10303);
nor NOR4 (N10308, N10287, N3204, N6236, N6881);
xor XOR2 (N10309, N10286, N5780);
buf BUF1 (N10310, N10280);
nand NAND4 (N10311, N10310, N7661, N8043, N9803);
xor XOR2 (N10312, N10300, N10171);
or OR4 (N10313, N10307, N7941, N7993, N5464);
nor NOR2 (N10314, N10299, N6176);
buf BUF1 (N10315, N10311);
not NOT1 (N10316, N10314);
buf BUF1 (N10317, N10309);
not NOT1 (N10318, N10306);
and AND4 (N10319, N10313, N7851, N2945, N1119);
or OR3 (N10320, N10298, N6172, N1834);
xor XOR2 (N10321, N10294, N7886);
nor NOR2 (N10322, N10320, N10291);
buf BUF1 (N10323, N10319);
nand NAND4 (N10324, N10321, N9313, N4938, N7166);
not NOT1 (N10325, N10317);
buf BUF1 (N10326, N10305);
and AND4 (N10327, N10323, N3371, N4923, N6658);
not NOT1 (N10328, N10318);
xor XOR2 (N10329, N10312, N5957);
and AND3 (N10330, N10329, N4687, N5754);
nor NOR3 (N10331, N10322, N2573, N8532);
not NOT1 (N10332, N10327);
not NOT1 (N10333, N10328);
buf BUF1 (N10334, N10308);
not NOT1 (N10335, N10326);
or OR2 (N10336, N10330, N2265);
buf BUF1 (N10337, N10335);
nand NAND2 (N10338, N10334, N1738);
or OR4 (N10339, N10316, N5307, N6644, N3644);
and AND3 (N10340, N10333, N8947, N2181);
not NOT1 (N10341, N10336);
or OR3 (N10342, N10338, N7048, N184);
nand NAND4 (N10343, N10337, N6592, N1431, N2001);
and AND3 (N10344, N10324, N2687, N8675);
xor XOR2 (N10345, N10325, N8090);
nor NOR4 (N10346, N10332, N8731, N10266, N9169);
or OR2 (N10347, N10342, N3994);
buf BUF1 (N10348, N10315);
buf BUF1 (N10349, N10345);
and AND3 (N10350, N10347, N524, N10239);
xor XOR2 (N10351, N10343, N3487);
and AND4 (N10352, N10344, N8113, N8612, N8952);
nor NOR3 (N10353, N10348, N6376, N7579);
xor XOR2 (N10354, N10351, N5993);
buf BUF1 (N10355, N10354);
nand NAND2 (N10356, N10350, N9159);
nand NAND3 (N10357, N10346, N376, N4646);
buf BUF1 (N10358, N10341);
nand NAND3 (N10359, N10353, N1877, N6338);
xor XOR2 (N10360, N10358, N5758);
xor XOR2 (N10361, N10339, N6455);
not NOT1 (N10362, N10361);
not NOT1 (N10363, N10340);
and AND4 (N10364, N10352, N6426, N1373, N10165);
xor XOR2 (N10365, N10355, N4057);
xor XOR2 (N10366, N10331, N3962);
nor NOR3 (N10367, N10363, N8692, N6701);
nor NOR3 (N10368, N10365, N9434, N9055);
nand NAND2 (N10369, N10360, N4615);
nand NAND3 (N10370, N10366, N8282, N3260);
not NOT1 (N10371, N10359);
nand NAND3 (N10372, N10369, N1376, N1583);
and AND2 (N10373, N10372, N1405);
nor NOR2 (N10374, N10356, N7318);
not NOT1 (N10375, N10368);
nand NAND2 (N10376, N10362, N5569);
not NOT1 (N10377, N10364);
nand NAND2 (N10378, N10375, N7961);
and AND3 (N10379, N10357, N710, N3212);
buf BUF1 (N10380, N10367);
buf BUF1 (N10381, N10373);
not NOT1 (N10382, N10376);
xor XOR2 (N10383, N10374, N3763);
buf BUF1 (N10384, N10378);
not NOT1 (N10385, N10381);
and AND4 (N10386, N10382, N1722, N9469, N2667);
buf BUF1 (N10387, N10377);
or OR3 (N10388, N10379, N2061, N2400);
or OR2 (N10389, N10388, N7009);
buf BUF1 (N10390, N10386);
or OR3 (N10391, N10385, N4531, N7505);
nand NAND3 (N10392, N10370, N5600, N7429);
nand NAND4 (N10393, N10391, N3437, N1375, N1759);
not NOT1 (N10394, N10392);
and AND3 (N10395, N10389, N9131, N4045);
nand NAND2 (N10396, N10349, N3972);
nor NOR4 (N10397, N10371, N6358, N5874, N3493);
nor NOR2 (N10398, N10397, N7018);
buf BUF1 (N10399, N10387);
xor XOR2 (N10400, N10380, N438);
not NOT1 (N10401, N10394);
or OR3 (N10402, N10393, N7339, N617);
not NOT1 (N10403, N10398);
nand NAND4 (N10404, N10396, N4746, N2142, N9374);
not NOT1 (N10405, N10383);
buf BUF1 (N10406, N10405);
nor NOR4 (N10407, N10401, N4626, N2367, N4747);
not NOT1 (N10408, N10384);
nand NAND4 (N10409, N10407, N3336, N7207, N3836);
nor NOR2 (N10410, N10402, N7943);
nor NOR2 (N10411, N10390, N8055);
xor XOR2 (N10412, N10399, N9275);
nand NAND4 (N10413, N10404, N3620, N4129, N2783);
or OR4 (N10414, N10400, N9740, N9660, N3478);
nand NAND2 (N10415, N10412, N1643);
buf BUF1 (N10416, N10408);
nor NOR2 (N10417, N10413, N3270);
and AND3 (N10418, N10414, N9570, N8090);
not NOT1 (N10419, N10411);
nor NOR4 (N10420, N10415, N9454, N2817, N8155);
buf BUF1 (N10421, N10419);
nor NOR3 (N10422, N10403, N9978, N3935);
or OR3 (N10423, N10409, N2780, N2952);
buf BUF1 (N10424, N10422);
or OR4 (N10425, N10423, N7577, N2588, N9439);
or OR2 (N10426, N10421, N7941);
xor XOR2 (N10427, N10420, N5363);
nand NAND3 (N10428, N10417, N3656, N7373);
or OR2 (N10429, N10428, N910);
xor XOR2 (N10430, N10410, N285);
not NOT1 (N10431, N10395);
nor NOR4 (N10432, N10427, N7321, N4371, N5271);
and AND2 (N10433, N10429, N535);
and AND3 (N10434, N10433, N8270, N10167);
not NOT1 (N10435, N10418);
or OR2 (N10436, N10426, N3616);
and AND4 (N10437, N10424, N482, N9846, N1688);
nand NAND2 (N10438, N10416, N5329);
buf BUF1 (N10439, N10434);
nand NAND3 (N10440, N10425, N5612, N7924);
xor XOR2 (N10441, N10406, N8924);
and AND2 (N10442, N10439, N9524);
nand NAND4 (N10443, N10436, N4163, N7478, N8078);
buf BUF1 (N10444, N10443);
or OR4 (N10445, N10444, N3250, N34, N4880);
or OR4 (N10446, N10432, N3488, N3587, N5953);
or OR2 (N10447, N10446, N4709);
and AND3 (N10448, N10438, N234, N8813);
and AND4 (N10449, N10437, N8738, N6742, N5507);
buf BUF1 (N10450, N10449);
and AND3 (N10451, N10445, N3746, N4206);
xor XOR2 (N10452, N10448, N7365);
or OR4 (N10453, N10452, N5564, N4615, N2521);
xor XOR2 (N10454, N10442, N7531);
nand NAND4 (N10455, N10435, N1310, N6857, N2417);
or OR2 (N10456, N10431, N1446);
nor NOR4 (N10457, N10430, N2278, N5681, N5831);
and AND4 (N10458, N10456, N3429, N10009, N204);
buf BUF1 (N10459, N10450);
nand NAND3 (N10460, N10447, N6345, N4473);
buf BUF1 (N10461, N10451);
xor XOR2 (N10462, N10457, N10190);
not NOT1 (N10463, N10453);
nor NOR2 (N10464, N10440, N936);
nand NAND3 (N10465, N10454, N1861, N6653);
or OR4 (N10466, N10465, N7887, N3982, N846);
xor XOR2 (N10467, N10441, N9615);
nand NAND2 (N10468, N10462, N1273);
buf BUF1 (N10469, N10459);
nand NAND2 (N10470, N10455, N5045);
buf BUF1 (N10471, N10470);
nand NAND4 (N10472, N10460, N3655, N1948, N4254);
buf BUF1 (N10473, N10466);
buf BUF1 (N10474, N10469);
xor XOR2 (N10475, N10471, N4886);
buf BUF1 (N10476, N10472);
nor NOR2 (N10477, N10461, N3816);
xor XOR2 (N10478, N10476, N8904);
buf BUF1 (N10479, N10474);
nand NAND3 (N10480, N10477, N110, N2664);
xor XOR2 (N10481, N10475, N10071);
nor NOR2 (N10482, N10463, N1784);
and AND4 (N10483, N10480, N3312, N8389, N1985);
xor XOR2 (N10484, N10458, N5550);
buf BUF1 (N10485, N10464);
xor XOR2 (N10486, N10479, N8722);
or OR3 (N10487, N10481, N3821, N3089);
xor XOR2 (N10488, N10478, N9488);
nand NAND3 (N10489, N10486, N10164, N6347);
nand NAND2 (N10490, N10473, N7831);
buf BUF1 (N10491, N10485);
buf BUF1 (N10492, N10484);
not NOT1 (N10493, N10483);
nand NAND2 (N10494, N10489, N9853);
and AND3 (N10495, N10468, N10173, N9549);
not NOT1 (N10496, N10467);
xor XOR2 (N10497, N10488, N5258);
nand NAND4 (N10498, N10495, N377, N1836, N6646);
not NOT1 (N10499, N10492);
and AND2 (N10500, N10487, N6772);
or OR4 (N10501, N10500, N4364, N9127, N1921);
not NOT1 (N10502, N10499);
nor NOR4 (N10503, N10493, N7203, N7011, N7552);
or OR2 (N10504, N10482, N7838);
not NOT1 (N10505, N10496);
not NOT1 (N10506, N10501);
and AND3 (N10507, N10497, N4886, N9646);
buf BUF1 (N10508, N10505);
or OR2 (N10509, N10506, N7026);
buf BUF1 (N10510, N10503);
nor NOR4 (N10511, N10502, N8092, N6521, N6487);
nor NOR2 (N10512, N10490, N2929);
not NOT1 (N10513, N10511);
nor NOR2 (N10514, N10491, N8680);
nand NAND3 (N10515, N10510, N8462, N1471);
buf BUF1 (N10516, N10494);
xor XOR2 (N10517, N10498, N6611);
and AND4 (N10518, N10514, N1004, N9645, N5177);
and AND3 (N10519, N10507, N4129, N4916);
or OR3 (N10520, N10518, N3790, N9263);
nor NOR4 (N10521, N10509, N5498, N5951, N10372);
or OR3 (N10522, N10517, N4634, N4408);
or OR2 (N10523, N10512, N760);
buf BUF1 (N10524, N10519);
nor NOR2 (N10525, N10523, N9371);
or OR4 (N10526, N10508, N716, N759, N8213);
nor NOR2 (N10527, N10515, N7796);
nor NOR4 (N10528, N10521, N5124, N8311, N8451);
xor XOR2 (N10529, N10527, N8214);
or OR4 (N10530, N10520, N10101, N576, N2847);
xor XOR2 (N10531, N10530, N3550);
buf BUF1 (N10532, N10529);
or OR2 (N10533, N10504, N9856);
xor XOR2 (N10534, N10528, N4856);
not NOT1 (N10535, N10526);
nand NAND3 (N10536, N10524, N4807, N2899);
xor XOR2 (N10537, N10532, N8748);
or OR3 (N10538, N10516, N8570, N5037);
nand NAND3 (N10539, N10513, N10254, N8694);
or OR3 (N10540, N10538, N5083, N6357);
not NOT1 (N10541, N10535);
nor NOR3 (N10542, N10522, N1470, N3271);
nor NOR3 (N10543, N10539, N8473, N6556);
xor XOR2 (N10544, N10525, N2073);
or OR3 (N10545, N10543, N8969, N1664);
not NOT1 (N10546, N10536);
xor XOR2 (N10547, N10541, N9259);
xor XOR2 (N10548, N10545, N5027);
xor XOR2 (N10549, N10542, N9323);
not NOT1 (N10550, N10531);
nor NOR2 (N10551, N10533, N3144);
xor XOR2 (N10552, N10537, N2964);
nor NOR3 (N10553, N10534, N2177, N6018);
buf BUF1 (N10554, N10550);
nor NOR2 (N10555, N10540, N4067);
not NOT1 (N10556, N10554);
not NOT1 (N10557, N10553);
and AND4 (N10558, N10549, N9365, N6983, N2769);
or OR2 (N10559, N10556, N8098);
nor NOR3 (N10560, N10547, N8037, N8172);
nand NAND3 (N10561, N10555, N9158, N3977);
xor XOR2 (N10562, N10546, N6594);
buf BUF1 (N10563, N10551);
or OR4 (N10564, N10563, N9519, N3273, N9230);
nor NOR2 (N10565, N10558, N7005);
nand NAND4 (N10566, N10559, N3393, N6713, N2776);
nor NOR2 (N10567, N10544, N3621);
xor XOR2 (N10568, N10564, N5185);
and AND4 (N10569, N10562, N3340, N6944, N7908);
buf BUF1 (N10570, N10561);
and AND4 (N10571, N10565, N5654, N4707, N9156);
nand NAND3 (N10572, N10567, N3730, N1287);
and AND3 (N10573, N10548, N2768, N3234);
and AND4 (N10574, N10573, N4560, N476, N6617);
and AND3 (N10575, N10571, N7692, N2209);
buf BUF1 (N10576, N10574);
or OR4 (N10577, N10560, N1447, N3586, N4109);
or OR3 (N10578, N10576, N442, N5144);
and AND2 (N10579, N10570, N10138);
xor XOR2 (N10580, N10566, N10374);
not NOT1 (N10581, N10552);
or OR4 (N10582, N10577, N5938, N6778, N8579);
and AND3 (N10583, N10582, N10153, N8565);
or OR3 (N10584, N10569, N4470, N2130);
nand NAND2 (N10585, N10583, N3180);
and AND2 (N10586, N10572, N3708);
and AND4 (N10587, N10585, N5124, N902, N7828);
buf BUF1 (N10588, N10579);
xor XOR2 (N10589, N10580, N4969);
nor NOR4 (N10590, N10578, N2841, N5687, N2584);
not NOT1 (N10591, N10584);
or OR3 (N10592, N10587, N1403, N8886);
and AND2 (N10593, N10586, N4325);
xor XOR2 (N10594, N10589, N5045);
not NOT1 (N10595, N10593);
not NOT1 (N10596, N10575);
and AND4 (N10597, N10591, N6041, N6636, N1610);
xor XOR2 (N10598, N10568, N1952);
xor XOR2 (N10599, N10581, N178);
not NOT1 (N10600, N10557);
and AND2 (N10601, N10599, N5512);
buf BUF1 (N10602, N10598);
xor XOR2 (N10603, N10590, N3598);
or OR4 (N10604, N10597, N3472, N8935, N5848);
not NOT1 (N10605, N10601);
xor XOR2 (N10606, N10600, N7908);
buf BUF1 (N10607, N10594);
nor NOR3 (N10608, N10595, N8273, N2294);
and AND4 (N10609, N10592, N757, N2066, N6449);
not NOT1 (N10610, N10603);
and AND4 (N10611, N10605, N7895, N5754, N7080);
nor NOR2 (N10612, N10588, N3925);
xor XOR2 (N10613, N10612, N3299);
xor XOR2 (N10614, N10604, N6171);
and AND2 (N10615, N10606, N307);
or OR4 (N10616, N10611, N7517, N9418, N2631);
nor NOR4 (N10617, N10596, N6523, N2768, N9084);
buf BUF1 (N10618, N10608);
nand NAND2 (N10619, N10615, N2696);
buf BUF1 (N10620, N10619);
xor XOR2 (N10621, N10602, N9730);
nor NOR3 (N10622, N10617, N7136, N6612);
not NOT1 (N10623, N10607);
buf BUF1 (N10624, N10610);
or OR4 (N10625, N10623, N9235, N6613, N10380);
or OR2 (N10626, N10613, N3348);
buf BUF1 (N10627, N10609);
and AND2 (N10628, N10625, N8135);
not NOT1 (N10629, N10628);
or OR3 (N10630, N10624, N960, N4684);
nor NOR3 (N10631, N10618, N8107, N7673);
buf BUF1 (N10632, N10621);
or OR3 (N10633, N10631, N742, N10429);
or OR2 (N10634, N10626, N7226);
xor XOR2 (N10635, N10616, N10558);
xor XOR2 (N10636, N10635, N7050);
or OR3 (N10637, N10622, N10240, N2954);
or OR4 (N10638, N10614, N3563, N4910, N10370);
not NOT1 (N10639, N10620);
nor NOR2 (N10640, N10636, N8539);
buf BUF1 (N10641, N10640);
not NOT1 (N10642, N10630);
not NOT1 (N10643, N10637);
buf BUF1 (N10644, N10629);
and AND2 (N10645, N10642, N5934);
and AND3 (N10646, N10634, N5372, N9949);
nand NAND4 (N10647, N10633, N339, N9743, N8834);
nand NAND3 (N10648, N10645, N4437, N9903);
nand NAND3 (N10649, N10632, N3799, N9834);
not NOT1 (N10650, N10644);
buf BUF1 (N10651, N10638);
and AND4 (N10652, N10649, N9708, N8555, N4666);
nor NOR4 (N10653, N10652, N9032, N9115, N1771);
xor XOR2 (N10654, N10653, N1360);
xor XOR2 (N10655, N10650, N8881);
not NOT1 (N10656, N10651);
xor XOR2 (N10657, N10656, N486);
nand NAND2 (N10658, N10655, N2249);
not NOT1 (N10659, N10658);
nand NAND2 (N10660, N10641, N1736);
xor XOR2 (N10661, N10648, N10476);
nor NOR3 (N10662, N10646, N4636, N2259);
xor XOR2 (N10663, N10654, N4958);
and AND2 (N10664, N10657, N4312);
nor NOR4 (N10665, N10647, N2694, N5938, N1444);
and AND2 (N10666, N10665, N7371);
not NOT1 (N10667, N10659);
not NOT1 (N10668, N10639);
or OR2 (N10669, N10666, N4417);
not NOT1 (N10670, N10627);
nor NOR3 (N10671, N10662, N4586, N9460);
not NOT1 (N10672, N10668);
buf BUF1 (N10673, N10667);
nor NOR4 (N10674, N10664, N10669, N1496, N2708);
xor XOR2 (N10675, N6301, N9242);
or OR3 (N10676, N10673, N4592, N2944);
or OR4 (N10677, N10643, N274, N7081, N8899);
not NOT1 (N10678, N10661);
buf BUF1 (N10679, N10660);
or OR3 (N10680, N10663, N124, N8686);
xor XOR2 (N10681, N10680, N6812);
nor NOR3 (N10682, N10672, N1195, N5836);
nand NAND3 (N10683, N10671, N10550, N3230);
and AND4 (N10684, N10675, N10181, N6076, N8784);
buf BUF1 (N10685, N10679);
buf BUF1 (N10686, N10685);
or OR2 (N10687, N10684, N5805);
nand NAND3 (N10688, N10687, N5880, N7283);
xor XOR2 (N10689, N10681, N3281);
or OR3 (N10690, N10678, N5666, N864);
xor XOR2 (N10691, N10674, N4505);
or OR2 (N10692, N10676, N8162);
nand NAND3 (N10693, N10677, N4421, N731);
not NOT1 (N10694, N10692);
nor NOR2 (N10695, N10689, N4165);
buf BUF1 (N10696, N10694);
buf BUF1 (N10697, N10690);
or OR4 (N10698, N10686, N6458, N9767, N8914);
and AND2 (N10699, N10682, N2079);
or OR4 (N10700, N10688, N8803, N3543, N7598);
and AND4 (N10701, N10691, N519, N352, N81);
and AND2 (N10702, N10701, N9280);
or OR3 (N10703, N10697, N5632, N7452);
and AND4 (N10704, N10698, N9155, N2098, N1606);
xor XOR2 (N10705, N10699, N1211);
nor NOR3 (N10706, N10693, N3627, N8507);
buf BUF1 (N10707, N10706);
and AND2 (N10708, N10670, N2956);
or OR4 (N10709, N10700, N10271, N9261, N4824);
not NOT1 (N10710, N10707);
not NOT1 (N10711, N10702);
nor NOR4 (N10712, N10696, N325, N1041, N686);
not NOT1 (N10713, N10705);
or OR4 (N10714, N10712, N5783, N2066, N2223);
and AND3 (N10715, N10703, N6287, N231);
not NOT1 (N10716, N10708);
buf BUF1 (N10717, N10715);
nand NAND3 (N10718, N10709, N1267, N4983);
nor NOR4 (N10719, N10718, N8900, N4128, N4213);
buf BUF1 (N10720, N10704);
buf BUF1 (N10721, N10720);
and AND4 (N10722, N10695, N3510, N8993, N6814);
xor XOR2 (N10723, N10710, N4807);
not NOT1 (N10724, N10713);
not NOT1 (N10725, N10721);
not NOT1 (N10726, N10714);
not NOT1 (N10727, N10726);
xor XOR2 (N10728, N10717, N7211);
nor NOR4 (N10729, N10723, N3491, N8037, N7071);
xor XOR2 (N10730, N10728, N1325);
or OR3 (N10731, N10729, N6982, N8764);
and AND3 (N10732, N10683, N668, N6406);
nor NOR4 (N10733, N10716, N3663, N3522, N3184);
nand NAND3 (N10734, N10733, N8824, N6150);
nor NOR4 (N10735, N10727, N8262, N2176, N5301);
not NOT1 (N10736, N10730);
nor NOR4 (N10737, N10736, N1180, N1540, N7424);
nor NOR3 (N10738, N10722, N4952, N516);
not NOT1 (N10739, N10732);
and AND4 (N10740, N10731, N7511, N7267, N2177);
nor NOR3 (N10741, N10719, N8035, N5381);
or OR2 (N10742, N10739, N9142);
or OR2 (N10743, N10711, N10661);
nor NOR3 (N10744, N10742, N3206, N2092);
xor XOR2 (N10745, N10737, N6217);
nor NOR3 (N10746, N10725, N8234, N2702);
xor XOR2 (N10747, N10738, N6403);
or OR3 (N10748, N10746, N10293, N7762);
nor NOR4 (N10749, N10734, N4651, N9913, N2425);
xor XOR2 (N10750, N10743, N10167);
buf BUF1 (N10751, N10740);
not NOT1 (N10752, N10751);
or OR4 (N10753, N10744, N4661, N2797, N5299);
not NOT1 (N10754, N10741);
and AND2 (N10755, N10750, N9684);
nand NAND4 (N10756, N10753, N9126, N6146, N8427);
xor XOR2 (N10757, N10735, N6642);
nand NAND2 (N10758, N10748, N6710);
not NOT1 (N10759, N10747);
not NOT1 (N10760, N10759);
and AND2 (N10761, N10756, N2456);
or OR3 (N10762, N10724, N7482, N9129);
xor XOR2 (N10763, N10762, N1694);
not NOT1 (N10764, N10763);
buf BUF1 (N10765, N10752);
not NOT1 (N10766, N10754);
not NOT1 (N10767, N10761);
nand NAND3 (N10768, N10764, N2304, N7516);
nand NAND3 (N10769, N10757, N3578, N1920);
buf BUF1 (N10770, N10766);
xor XOR2 (N10771, N10767, N2321);
buf BUF1 (N10772, N10765);
nand NAND2 (N10773, N10768, N5960);
nand NAND3 (N10774, N10760, N297, N612);
nor NOR4 (N10775, N10774, N8697, N10084, N3577);
nor NOR4 (N10776, N10769, N8798, N373, N1185);
or OR4 (N10777, N10770, N9553, N1980, N7921);
not NOT1 (N10778, N10772);
buf BUF1 (N10779, N10758);
not NOT1 (N10780, N10771);
nand NAND4 (N10781, N10778, N1998, N2318, N5858);
buf BUF1 (N10782, N10755);
nand NAND2 (N10783, N10775, N7143);
buf BUF1 (N10784, N10773);
nand NAND4 (N10785, N10777, N6595, N6381, N3751);
buf BUF1 (N10786, N10781);
nor NOR3 (N10787, N10745, N1884, N6617);
and AND4 (N10788, N10782, N1031, N758, N5368);
or OR2 (N10789, N10788, N8371);
nand NAND3 (N10790, N10779, N2100, N5329);
nor NOR4 (N10791, N10786, N4335, N9039, N6653);
nand NAND2 (N10792, N10790, N7709);
xor XOR2 (N10793, N10776, N1885);
xor XOR2 (N10794, N10792, N4527);
not NOT1 (N10795, N10789);
nand NAND2 (N10796, N10784, N7316);
buf BUF1 (N10797, N10785);
and AND2 (N10798, N10780, N4355);
or OR2 (N10799, N10794, N7604);
and AND2 (N10800, N10799, N5405);
buf BUF1 (N10801, N10800);
xor XOR2 (N10802, N10795, N5902);
nand NAND4 (N10803, N10798, N6703, N8612, N10651);
nor NOR2 (N10804, N10787, N8900);
or OR2 (N10805, N10797, N3082);
or OR4 (N10806, N10796, N1542, N2127, N3178);
nand NAND2 (N10807, N10805, N3761);
nand NAND3 (N10808, N10802, N2571, N3422);
nand NAND2 (N10809, N10791, N248);
buf BUF1 (N10810, N10804);
not NOT1 (N10811, N10783);
nand NAND3 (N10812, N10806, N4915, N3782);
nand NAND3 (N10813, N10811, N837, N7360);
or OR3 (N10814, N10749, N2579, N6486);
not NOT1 (N10815, N10809);
or OR4 (N10816, N10815, N10310, N6852, N6831);
and AND4 (N10817, N10813, N8406, N922, N10148);
nand NAND3 (N10818, N10807, N2428, N7620);
nand NAND4 (N10819, N10801, N3790, N9329, N4560);
xor XOR2 (N10820, N10817, N3085);
nand NAND2 (N10821, N10820, N4418);
xor XOR2 (N10822, N10808, N4174);
buf BUF1 (N10823, N10816);
xor XOR2 (N10824, N10823, N6175);
nand NAND3 (N10825, N10814, N1493, N8070);
or OR4 (N10826, N10812, N7191, N8117, N10614);
nand NAND2 (N10827, N10822, N7242);
nand NAND2 (N10828, N10819, N6597);
nand NAND4 (N10829, N10826, N7819, N1989, N442);
nand NAND3 (N10830, N10827, N3420, N5466);
buf BUF1 (N10831, N10829);
or OR4 (N10832, N10830, N3667, N881, N6449);
not NOT1 (N10833, N10825);
not NOT1 (N10834, N10793);
xor XOR2 (N10835, N10833, N662);
nand NAND4 (N10836, N10832, N6173, N7747, N8909);
or OR3 (N10837, N10824, N10214, N8898);
and AND2 (N10838, N10831, N6360);
or OR3 (N10839, N10828, N7905, N3117);
nand NAND2 (N10840, N10838, N7592);
and AND3 (N10841, N10810, N2806, N3437);
and AND4 (N10842, N10836, N5865, N10265, N9335);
nor NOR3 (N10843, N10842, N7693, N1519);
buf BUF1 (N10844, N10818);
nor NOR2 (N10845, N10839, N8399);
and AND3 (N10846, N10834, N9150, N3220);
nor NOR3 (N10847, N10837, N5170, N2897);
and AND2 (N10848, N10821, N3816);
not NOT1 (N10849, N10840);
nor NOR4 (N10850, N10803, N543, N4188, N10004);
and AND4 (N10851, N10849, N7599, N2119, N6203);
buf BUF1 (N10852, N10846);
buf BUF1 (N10853, N10848);
or OR4 (N10854, N10850, N4952, N2913, N2328);
not NOT1 (N10855, N10851);
not NOT1 (N10856, N10845);
not NOT1 (N10857, N10852);
or OR2 (N10858, N10841, N9706);
or OR3 (N10859, N10844, N840, N8803);
xor XOR2 (N10860, N10843, N3245);
buf BUF1 (N10861, N10858);
and AND3 (N10862, N10853, N1265, N2432);
buf BUF1 (N10863, N10847);
nand NAND4 (N10864, N10859, N4547, N1820, N9714);
xor XOR2 (N10865, N10835, N4221);
or OR3 (N10866, N10864, N975, N9848);
and AND4 (N10867, N10857, N4874, N10365, N1229);
not NOT1 (N10868, N10861);
nand NAND3 (N10869, N10867, N2043, N5223);
buf BUF1 (N10870, N10865);
and AND3 (N10871, N10856, N8747, N7830);
nand NAND4 (N10872, N10870, N6382, N7261, N2943);
or OR2 (N10873, N10862, N5116);
and AND2 (N10874, N10868, N3629);
xor XOR2 (N10875, N10873, N9232);
or OR3 (N10876, N10874, N4270, N3598);
nand NAND4 (N10877, N10869, N8581, N8911, N3621);
buf BUF1 (N10878, N10866);
not NOT1 (N10879, N10876);
xor XOR2 (N10880, N10855, N64);
nor NOR2 (N10881, N10854, N9080);
not NOT1 (N10882, N10881);
nor NOR2 (N10883, N10871, N4351);
xor XOR2 (N10884, N10878, N8740);
buf BUF1 (N10885, N10872);
nor NOR2 (N10886, N10860, N5306);
nor NOR2 (N10887, N10885, N564);
nand NAND2 (N10888, N10887, N7280);
buf BUF1 (N10889, N10879);
and AND3 (N10890, N10877, N5809, N8265);
or OR4 (N10891, N10888, N9220, N9417, N8232);
and AND2 (N10892, N10886, N5768);
nand NAND3 (N10893, N10884, N6628, N5968);
buf BUF1 (N10894, N10892);
or OR2 (N10895, N10875, N8018);
not NOT1 (N10896, N10882);
and AND3 (N10897, N10889, N10143, N3516);
and AND4 (N10898, N10863, N4733, N7754, N6521);
nand NAND2 (N10899, N10883, N2695);
buf BUF1 (N10900, N10891);
buf BUF1 (N10901, N10898);
xor XOR2 (N10902, N10894, N1057);
or OR3 (N10903, N10895, N6561, N2286);
not NOT1 (N10904, N10901);
nor NOR4 (N10905, N10899, N871, N10511, N10347);
buf BUF1 (N10906, N10902);
nand NAND3 (N10907, N10893, N5242, N7715);
xor XOR2 (N10908, N10903, N4199);
xor XOR2 (N10909, N10907, N343);
not NOT1 (N10910, N10896);
nor NOR4 (N10911, N10908, N3970, N1219, N4064);
buf BUF1 (N10912, N10905);
nand NAND2 (N10913, N10909, N8183);
not NOT1 (N10914, N10912);
or OR4 (N10915, N10910, N6822, N6354, N9615);
not NOT1 (N10916, N10913);
or OR2 (N10917, N10900, N2448);
nand NAND4 (N10918, N10915, N5545, N798, N5349);
nor NOR2 (N10919, N10890, N3338);
nand NAND4 (N10920, N10918, N2324, N9178, N9962);
or OR3 (N10921, N10880, N8382, N4939);
or OR2 (N10922, N10906, N2203);
not NOT1 (N10923, N10897);
nor NOR3 (N10924, N10920, N9128, N6075);
nor NOR2 (N10925, N10923, N5642);
nand NAND2 (N10926, N10925, N9934);
nor NOR4 (N10927, N10916, N5030, N10636, N8097);
and AND4 (N10928, N10919, N5993, N4602, N2331);
not NOT1 (N10929, N10917);
or OR2 (N10930, N10926, N252);
and AND3 (N10931, N10911, N2069, N1076);
xor XOR2 (N10932, N10930, N7206);
buf BUF1 (N10933, N10914);
or OR3 (N10934, N10932, N10004, N5581);
buf BUF1 (N10935, N10934);
nand NAND3 (N10936, N10935, N720, N8032);
or OR3 (N10937, N10936, N9493, N396);
nand NAND2 (N10938, N10937, N7303);
or OR2 (N10939, N10904, N3492);
nor NOR4 (N10940, N10924, N4736, N1861, N6462);
xor XOR2 (N10941, N10931, N1005);
nor NOR4 (N10942, N10938, N4508, N4218, N7307);
xor XOR2 (N10943, N10928, N4243);
or OR3 (N10944, N10942, N10593, N9505);
nor NOR3 (N10945, N10927, N9954, N5055);
xor XOR2 (N10946, N10944, N6216);
nand NAND2 (N10947, N10941, N3298);
buf BUF1 (N10948, N10945);
buf BUF1 (N10949, N10933);
nor NOR3 (N10950, N10948, N4119, N5979);
xor XOR2 (N10951, N10946, N472);
or OR4 (N10952, N10943, N8500, N9136, N5244);
and AND2 (N10953, N10951, N4514);
not NOT1 (N10954, N10940);
and AND4 (N10955, N10922, N3680, N5176, N2129);
or OR4 (N10956, N10921, N9672, N6448, N2317);
nand NAND3 (N10957, N10950, N7800, N4700);
and AND2 (N10958, N10929, N8523);
buf BUF1 (N10959, N10957);
xor XOR2 (N10960, N10955, N4823);
not NOT1 (N10961, N10953);
buf BUF1 (N10962, N10956);
not NOT1 (N10963, N10959);
nor NOR4 (N10964, N10952, N5574, N8068, N1616);
not NOT1 (N10965, N10960);
not NOT1 (N10966, N10949);
xor XOR2 (N10967, N10961, N8202);
not NOT1 (N10968, N10962);
or OR3 (N10969, N10939, N8349, N6891);
and AND2 (N10970, N10958, N1647);
and AND2 (N10971, N10968, N5864);
nand NAND2 (N10972, N10963, N6792);
buf BUF1 (N10973, N10954);
buf BUF1 (N10974, N10973);
buf BUF1 (N10975, N10974);
not NOT1 (N10976, N10947);
nor NOR4 (N10977, N10972, N4447, N8031, N2557);
xor XOR2 (N10978, N10971, N4779);
nor NOR2 (N10979, N10969, N8092);
or OR2 (N10980, N10979, N969);
nor NOR4 (N10981, N10980, N4407, N4380, N4909);
buf BUF1 (N10982, N10977);
buf BUF1 (N10983, N10978);
buf BUF1 (N10984, N10975);
not NOT1 (N10985, N10966);
or OR2 (N10986, N10983, N9056);
xor XOR2 (N10987, N10986, N5644);
buf BUF1 (N10988, N10982);
xor XOR2 (N10989, N10964, N10806);
nand NAND3 (N10990, N10988, N8174, N4033);
and AND3 (N10991, N10976, N419, N7582);
nor NOR2 (N10992, N10970, N1705);
nor NOR4 (N10993, N10990, N7968, N9564, N5549);
and AND4 (N10994, N10967, N7669, N1658, N7098);
nand NAND3 (N10995, N10991, N4494, N1975);
buf BUF1 (N10996, N10987);
or OR3 (N10997, N10981, N4872, N6902);
xor XOR2 (N10998, N10995, N7282);
nand NAND2 (N10999, N10996, N849);
xor XOR2 (N11000, N10998, N2904);
nor NOR2 (N11001, N11000, N3628);
not NOT1 (N11002, N10989);
or OR3 (N11003, N10999, N10204, N519);
buf BUF1 (N11004, N10992);
buf BUF1 (N11005, N10994);
xor XOR2 (N11006, N11005, N4749);
nor NOR4 (N11007, N11001, N4877, N5477, N7034);
nand NAND2 (N11008, N10997, N4400);
and AND3 (N11009, N11008, N9755, N2610);
not NOT1 (N11010, N11004);
or OR2 (N11011, N11009, N9956);
nor NOR4 (N11012, N11007, N4344, N289, N4321);
buf BUF1 (N11013, N10984);
nor NOR4 (N11014, N11006, N9939, N7054, N1430);
not NOT1 (N11015, N11011);
nand NAND3 (N11016, N10993, N89, N2569);
buf BUF1 (N11017, N11012);
not NOT1 (N11018, N11002);
nand NAND2 (N11019, N11014, N8102);
xor XOR2 (N11020, N10965, N7552);
not NOT1 (N11021, N11019);
or OR3 (N11022, N11021, N10992, N6255);
or OR4 (N11023, N11020, N9921, N10158, N6097);
not NOT1 (N11024, N11003);
buf BUF1 (N11025, N10985);
not NOT1 (N11026, N11015);
not NOT1 (N11027, N11017);
buf BUF1 (N11028, N11018);
xor XOR2 (N11029, N11022, N7038);
xor XOR2 (N11030, N11029, N10964);
or OR2 (N11031, N11024, N3008);
nor NOR4 (N11032, N11026, N9421, N8137, N9763);
buf BUF1 (N11033, N11030);
or OR4 (N11034, N11028, N4034, N6822, N3578);
or OR3 (N11035, N11031, N8340, N1151);
and AND4 (N11036, N11023, N6490, N445, N5973);
xor XOR2 (N11037, N11034, N10650);
buf BUF1 (N11038, N11010);
nor NOR4 (N11039, N11027, N5153, N6855, N10768);
nand NAND4 (N11040, N11037, N7756, N5574, N3068);
and AND4 (N11041, N11040, N6540, N61, N7778);
xor XOR2 (N11042, N11035, N4247);
or OR3 (N11043, N11042, N1241, N6492);
nor NOR2 (N11044, N11041, N7894);
xor XOR2 (N11045, N11038, N9283);
or OR4 (N11046, N11045, N9470, N3242, N6924);
or OR2 (N11047, N11046, N9133);
or OR3 (N11048, N11036, N68, N2830);
or OR4 (N11049, N11044, N7918, N7479, N5327);
and AND3 (N11050, N11033, N8125, N8677);
nand NAND2 (N11051, N11049, N3177);
not NOT1 (N11052, N11047);
nor NOR3 (N11053, N11043, N3385, N725);
nor NOR2 (N11054, N11013, N9344);
not NOT1 (N11055, N11051);
and AND3 (N11056, N11053, N4798, N10406);
nand NAND4 (N11057, N11052, N6840, N9274, N3366);
xor XOR2 (N11058, N11056, N6840);
and AND4 (N11059, N11055, N1824, N322, N9637);
or OR2 (N11060, N11048, N6915);
or OR3 (N11061, N11058, N8022, N2417);
xor XOR2 (N11062, N11039, N10020);
or OR3 (N11063, N11025, N1280, N3501);
not NOT1 (N11064, N11032);
xor XOR2 (N11065, N11062, N2934);
nor NOR4 (N11066, N11065, N4855, N2213, N9130);
nor NOR2 (N11067, N11060, N7815);
not NOT1 (N11068, N11054);
and AND3 (N11069, N11064, N1018, N3745);
xor XOR2 (N11070, N11050, N4520);
nor NOR4 (N11071, N11059, N792, N4486, N9622);
nand NAND2 (N11072, N11067, N3961);
buf BUF1 (N11073, N11072);
not NOT1 (N11074, N11063);
and AND3 (N11075, N11066, N7305, N2628);
buf BUF1 (N11076, N11075);
xor XOR2 (N11077, N11070, N7192);
xor XOR2 (N11078, N11068, N10898);
buf BUF1 (N11079, N11077);
buf BUF1 (N11080, N11069);
or OR3 (N11081, N11080, N8098, N6199);
nand NAND2 (N11082, N11061, N10798);
nor NOR3 (N11083, N11071, N6967, N1710);
or OR3 (N11084, N11079, N5824, N5801);
xor XOR2 (N11085, N11084, N837);
not NOT1 (N11086, N11057);
nor NOR3 (N11087, N11085, N1990, N934);
xor XOR2 (N11088, N11076, N3837);
or OR3 (N11089, N11082, N9412, N10602);
and AND4 (N11090, N11078, N1746, N6853, N9501);
and AND3 (N11091, N11090, N8072, N11090);
not NOT1 (N11092, N11089);
nand NAND2 (N11093, N11092, N1236);
or OR4 (N11094, N11016, N8264, N10147, N3116);
xor XOR2 (N11095, N11086, N9992);
nor NOR3 (N11096, N11087, N7122, N8539);
xor XOR2 (N11097, N11091, N6405);
nand NAND4 (N11098, N11081, N3463, N8452, N5935);
buf BUF1 (N11099, N11093);
xor XOR2 (N11100, N11074, N9460);
buf BUF1 (N11101, N11095);
nand NAND2 (N11102, N11101, N10988);
buf BUF1 (N11103, N11099);
buf BUF1 (N11104, N11097);
buf BUF1 (N11105, N11073);
nand NAND4 (N11106, N11100, N4638, N6959, N3336);
or OR4 (N11107, N11096, N5539, N1568, N6746);
nor NOR4 (N11108, N11102, N6887, N10008, N10887);
nand NAND2 (N11109, N11094, N1504);
nand NAND4 (N11110, N11105, N1596, N7209, N5235);
not NOT1 (N11111, N11109);
nand NAND2 (N11112, N11110, N2414);
or OR4 (N11113, N11103, N1682, N4681, N5454);
not NOT1 (N11114, N11112);
and AND2 (N11115, N11083, N8662);
and AND2 (N11116, N11106, N4578);
not NOT1 (N11117, N11098);
buf BUF1 (N11118, N11115);
nand NAND2 (N11119, N11114, N6901);
and AND2 (N11120, N11116, N3251);
or OR2 (N11121, N11113, N4652);
buf BUF1 (N11122, N11119);
xor XOR2 (N11123, N11118, N2979);
not NOT1 (N11124, N11117);
not NOT1 (N11125, N11108);
nand NAND3 (N11126, N11088, N2265, N10527);
nand NAND3 (N11127, N11121, N1212, N4994);
buf BUF1 (N11128, N11111);
not NOT1 (N11129, N11124);
buf BUF1 (N11130, N11120);
xor XOR2 (N11131, N11104, N8152);
or OR2 (N11132, N11107, N3959);
or OR2 (N11133, N11126, N1372);
nand NAND4 (N11134, N11131, N3226, N7923, N10402);
not NOT1 (N11135, N11125);
nand NAND2 (N11136, N11129, N5116);
nor NOR2 (N11137, N11135, N8541);
buf BUF1 (N11138, N11127);
not NOT1 (N11139, N11136);
xor XOR2 (N11140, N11138, N1332);
xor XOR2 (N11141, N11140, N7197);
nand NAND4 (N11142, N11134, N6226, N4094, N10887);
buf BUF1 (N11143, N11122);
nor NOR4 (N11144, N11139, N1863, N579, N10968);
or OR2 (N11145, N11128, N3604);
nand NAND2 (N11146, N11145, N9829);
and AND2 (N11147, N11133, N5450);
nor NOR2 (N11148, N11141, N3534);
and AND2 (N11149, N11144, N7156);
buf BUF1 (N11150, N11149);
not NOT1 (N11151, N11123);
or OR2 (N11152, N11147, N823);
and AND2 (N11153, N11130, N2153);
buf BUF1 (N11154, N11151);
nor NOR2 (N11155, N11150, N10510);
nand NAND2 (N11156, N11148, N1581);
nand NAND4 (N11157, N11152, N4005, N5766, N3570);
nand NAND2 (N11158, N11146, N6934);
buf BUF1 (N11159, N11132);
not NOT1 (N11160, N11142);
nand NAND2 (N11161, N11137, N4307);
nor NOR2 (N11162, N11155, N913);
or OR4 (N11163, N11159, N1348, N3066, N363);
and AND2 (N11164, N11163, N10599);
or OR2 (N11165, N11161, N2292);
and AND4 (N11166, N11164, N8171, N2673, N536);
and AND3 (N11167, N11143, N333, N6249);
or OR2 (N11168, N11160, N8720);
nor NOR2 (N11169, N11158, N6011);
xor XOR2 (N11170, N11154, N6786);
and AND3 (N11171, N11168, N1186, N6312);
nor NOR2 (N11172, N11171, N9888);
and AND4 (N11173, N11157, N5646, N3196, N1486);
nor NOR4 (N11174, N11153, N9046, N2817, N5865);
nand NAND3 (N11175, N11170, N7898, N5080);
or OR3 (N11176, N11167, N5905, N1675);
and AND2 (N11177, N11174, N2265);
not NOT1 (N11178, N11172);
xor XOR2 (N11179, N11169, N561);
xor XOR2 (N11180, N11173, N1369);
and AND3 (N11181, N11176, N11156, N3976);
nand NAND3 (N11182, N9596, N11024, N7635);
xor XOR2 (N11183, N11177, N10490);
nand NAND4 (N11184, N11166, N2583, N2511, N3312);
xor XOR2 (N11185, N11175, N6968);
nand NAND4 (N11186, N11184, N8153, N3335, N5277);
not NOT1 (N11187, N11165);
nand NAND4 (N11188, N11182, N3335, N3036, N7586);
and AND3 (N11189, N11162, N9199, N9989);
not NOT1 (N11190, N11183);
buf BUF1 (N11191, N11187);
nand NAND3 (N11192, N11186, N5246, N6614);
and AND4 (N11193, N11181, N48, N8280, N9236);
nor NOR2 (N11194, N11179, N7586);
and AND4 (N11195, N11193, N6518, N1025, N8788);
nor NOR2 (N11196, N11190, N8679);
xor XOR2 (N11197, N11196, N2194);
or OR4 (N11198, N11189, N2118, N1587, N7111);
not NOT1 (N11199, N11194);
or OR4 (N11200, N11185, N3439, N5870, N7900);
nor NOR2 (N11201, N11178, N11181);
and AND3 (N11202, N11195, N4648, N6707);
nor NOR3 (N11203, N11200, N10529, N1001);
nand NAND4 (N11204, N11199, N2203, N2725, N2586);
nand NAND4 (N11205, N11198, N5771, N7369, N3874);
not NOT1 (N11206, N11203);
nor NOR4 (N11207, N11202, N7042, N2903, N2375);
nor NOR4 (N11208, N11206, N2431, N2944, N6413);
or OR4 (N11209, N11191, N9376, N2176, N3644);
xor XOR2 (N11210, N11209, N4554);
and AND3 (N11211, N11207, N4605, N5210);
xor XOR2 (N11212, N11180, N8668);
or OR3 (N11213, N11204, N3084, N1097);
nand NAND2 (N11214, N11212, N6152);
nor NOR2 (N11215, N11214, N4344);
and AND3 (N11216, N11201, N6840, N61);
nand NAND4 (N11217, N11213, N4890, N6258, N1305);
nand NAND3 (N11218, N11197, N7338, N6190);
nand NAND2 (N11219, N11215, N2401);
or OR2 (N11220, N11216, N1741);
not NOT1 (N11221, N11192);
buf BUF1 (N11222, N11210);
and AND4 (N11223, N11218, N7952, N9749, N113);
nand NAND4 (N11224, N11219, N8002, N3023, N10828);
buf BUF1 (N11225, N11211);
and AND2 (N11226, N11225, N4);
or OR4 (N11227, N11208, N9997, N10090, N10486);
xor XOR2 (N11228, N11224, N7790);
not NOT1 (N11229, N11205);
xor XOR2 (N11230, N11221, N1470);
nand NAND3 (N11231, N11223, N10133, N8127);
nand NAND4 (N11232, N11229, N3187, N4368, N5532);
nand NAND2 (N11233, N11231, N508);
or OR4 (N11234, N11227, N8989, N1846, N6345);
nor NOR4 (N11235, N11217, N7749, N9307, N10598);
nand NAND4 (N11236, N11222, N1066, N1240, N8287);
nor NOR2 (N11237, N11232, N1048);
nor NOR4 (N11238, N11188, N4898, N10317, N2177);
buf BUF1 (N11239, N11228);
nor NOR3 (N11240, N11220, N5133, N1343);
buf BUF1 (N11241, N11239);
nand NAND4 (N11242, N11237, N8015, N10634, N4256);
xor XOR2 (N11243, N11242, N6942);
and AND2 (N11244, N11236, N6998);
nor NOR4 (N11245, N11241, N5019, N3292, N6483);
or OR2 (N11246, N11235, N7483);
not NOT1 (N11247, N11234);
xor XOR2 (N11248, N11238, N10879);
or OR2 (N11249, N11226, N4658);
nor NOR3 (N11250, N11248, N8627, N8117);
nor NOR2 (N11251, N11245, N824);
not NOT1 (N11252, N11249);
buf BUF1 (N11253, N11251);
nor NOR2 (N11254, N11240, N4774);
or OR4 (N11255, N11246, N9157, N6018, N3044);
and AND2 (N11256, N11253, N10501);
or OR2 (N11257, N11250, N6852);
not NOT1 (N11258, N11256);
nand NAND3 (N11259, N11244, N8011, N9606);
or OR2 (N11260, N11259, N408);
not NOT1 (N11261, N11233);
nand NAND3 (N11262, N11258, N9734, N10353);
xor XOR2 (N11263, N11261, N4448);
nor NOR4 (N11264, N11252, N4003, N42, N9057);
xor XOR2 (N11265, N11243, N4442);
or OR4 (N11266, N11262, N9168, N11252, N6751);
and AND2 (N11267, N11266, N1197);
buf BUF1 (N11268, N11257);
buf BUF1 (N11269, N11264);
buf BUF1 (N11270, N11254);
nor NOR4 (N11271, N11267, N9655, N11223, N9526);
xor XOR2 (N11272, N11230, N2352);
xor XOR2 (N11273, N11268, N4223);
or OR3 (N11274, N11263, N8072, N2138);
not NOT1 (N11275, N11247);
nand NAND2 (N11276, N11273, N3862);
or OR4 (N11277, N11260, N425, N3724, N11052);
xor XOR2 (N11278, N11275, N6506);
buf BUF1 (N11279, N11271);
not NOT1 (N11280, N11274);
or OR3 (N11281, N11270, N6912, N785);
nor NOR3 (N11282, N11276, N893, N2413);
nor NOR3 (N11283, N11279, N8508, N11232);
and AND3 (N11284, N11277, N6624, N6737);
and AND3 (N11285, N11284, N3483, N8105);
nand NAND4 (N11286, N11269, N2364, N1500, N6278);
not NOT1 (N11287, N11255);
not NOT1 (N11288, N11282);
nand NAND4 (N11289, N11278, N6833, N9371, N7457);
buf BUF1 (N11290, N11287);
xor XOR2 (N11291, N11289, N8545);
or OR4 (N11292, N11291, N1171, N10755, N4821);
or OR2 (N11293, N11288, N8442);
xor XOR2 (N11294, N11281, N5743);
or OR3 (N11295, N11286, N10802, N1214);
not NOT1 (N11296, N11290);
nand NAND4 (N11297, N11272, N9371, N3798, N3220);
buf BUF1 (N11298, N11293);
or OR4 (N11299, N11296, N3965, N1464, N5840);
xor XOR2 (N11300, N11294, N6553);
not NOT1 (N11301, N11285);
xor XOR2 (N11302, N11300, N7927);
buf BUF1 (N11303, N11283);
not NOT1 (N11304, N11302);
xor XOR2 (N11305, N11301, N9712);
nor NOR2 (N11306, N11295, N7934);
xor XOR2 (N11307, N11298, N6956);
nor NOR4 (N11308, N11265, N6266, N7834, N6456);
or OR3 (N11309, N11307, N11192, N5173);
nor NOR3 (N11310, N11292, N7825, N8186);
xor XOR2 (N11311, N11306, N338);
and AND3 (N11312, N11297, N6232, N5468);
nor NOR2 (N11313, N11309, N372);
or OR3 (N11314, N11312, N4928, N8765);
or OR4 (N11315, N11310, N7570, N1836, N879);
nor NOR2 (N11316, N11280, N7580);
nand NAND4 (N11317, N11299, N5799, N5800, N5216);
nand NAND3 (N11318, N11314, N3140, N10943);
xor XOR2 (N11319, N11318, N1865);
not NOT1 (N11320, N11316);
xor XOR2 (N11321, N11319, N5588);
xor XOR2 (N11322, N11308, N6639);
nor NOR4 (N11323, N11322, N4457, N5625, N8446);
nand NAND3 (N11324, N11315, N1181, N11079);
nand NAND2 (N11325, N11303, N7898);
not NOT1 (N11326, N11317);
or OR4 (N11327, N11323, N10098, N7767, N8104);
buf BUF1 (N11328, N11324);
xor XOR2 (N11329, N11311, N3429);
nand NAND2 (N11330, N11320, N4191);
and AND2 (N11331, N11321, N4444);
and AND3 (N11332, N11325, N6826, N4796);
not NOT1 (N11333, N11327);
nand NAND2 (N11334, N11332, N8186);
nand NAND3 (N11335, N11328, N2326, N8577);
nand NAND3 (N11336, N11326, N4185, N7866);
xor XOR2 (N11337, N11305, N3173);
nand NAND4 (N11338, N11331, N8256, N5370, N11241);
nand NAND3 (N11339, N11329, N10975, N1283);
nor NOR4 (N11340, N11313, N6860, N9175, N4382);
not NOT1 (N11341, N11337);
or OR2 (N11342, N11304, N1130);
xor XOR2 (N11343, N11334, N8436);
nand NAND4 (N11344, N11341, N9819, N9798, N6910);
or OR4 (N11345, N11336, N10609, N756, N8103);
nor NOR4 (N11346, N11340, N10259, N1761, N9898);
xor XOR2 (N11347, N11335, N439);
xor XOR2 (N11348, N11346, N2298);
and AND4 (N11349, N11344, N650, N483, N9106);
not NOT1 (N11350, N11338);
buf BUF1 (N11351, N11343);
xor XOR2 (N11352, N11342, N5899);
buf BUF1 (N11353, N11330);
nand NAND4 (N11354, N11349, N4830, N9114, N9156);
not NOT1 (N11355, N11351);
xor XOR2 (N11356, N11355, N9985);
or OR3 (N11357, N11356, N1752, N10451);
or OR4 (N11358, N11352, N5409, N2131, N8129);
xor XOR2 (N11359, N11350, N2291);
nor NOR4 (N11360, N11357, N9998, N665, N8934);
nand NAND4 (N11361, N11345, N10427, N3452, N2991);
xor XOR2 (N11362, N11360, N3326);
not NOT1 (N11363, N11353);
xor XOR2 (N11364, N11359, N4715);
nor NOR2 (N11365, N11358, N9283);
nor NOR4 (N11366, N11347, N4090, N2151, N10222);
buf BUF1 (N11367, N11333);
or OR3 (N11368, N11354, N8604, N7584);
nor NOR4 (N11369, N11367, N10656, N6068, N9701);
xor XOR2 (N11370, N11364, N4798);
xor XOR2 (N11371, N11366, N3285);
xor XOR2 (N11372, N11371, N5592);
buf BUF1 (N11373, N11363);
nor NOR3 (N11374, N11370, N5358, N5110);
and AND4 (N11375, N11365, N4966, N3055, N128);
nand NAND4 (N11376, N11361, N3733, N10436, N6436);
buf BUF1 (N11377, N11373);
or OR4 (N11378, N11348, N7210, N2822, N4358);
buf BUF1 (N11379, N11339);
xor XOR2 (N11380, N11374, N2371);
nand NAND2 (N11381, N11369, N9050);
xor XOR2 (N11382, N11372, N5765);
nor NOR3 (N11383, N11380, N4555, N5490);
not NOT1 (N11384, N11383);
nor NOR2 (N11385, N11376, N3138);
buf BUF1 (N11386, N11384);
or OR2 (N11387, N11368, N11226);
nand NAND3 (N11388, N11387, N6495, N1212);
nor NOR2 (N11389, N11377, N2915);
buf BUF1 (N11390, N11386);
or OR2 (N11391, N11390, N9769);
not NOT1 (N11392, N11389);
and AND3 (N11393, N11378, N5269, N4677);
and AND4 (N11394, N11391, N10570, N4017, N8678);
or OR4 (N11395, N11388, N7826, N4296, N121);
or OR3 (N11396, N11362, N951, N3587);
buf BUF1 (N11397, N11385);
and AND2 (N11398, N11395, N5265);
or OR4 (N11399, N11381, N1869, N10162, N4988);
and AND3 (N11400, N11393, N2033, N5903);
not NOT1 (N11401, N11396);
not NOT1 (N11402, N11394);
buf BUF1 (N11403, N11401);
or OR2 (N11404, N11400, N1613);
xor XOR2 (N11405, N11397, N4072);
or OR2 (N11406, N11402, N788);
xor XOR2 (N11407, N11406, N3841);
or OR2 (N11408, N11375, N1525);
or OR2 (N11409, N11404, N8756);
and AND2 (N11410, N11399, N10436);
xor XOR2 (N11411, N11379, N1618);
buf BUF1 (N11412, N11408);
or OR4 (N11413, N11407, N6432, N3742, N10514);
not NOT1 (N11414, N11405);
and AND3 (N11415, N11409, N9986, N1497);
buf BUF1 (N11416, N11398);
xor XOR2 (N11417, N11411, N1422);
xor XOR2 (N11418, N11392, N276);
nor NOR3 (N11419, N11416, N725, N2486);
not NOT1 (N11420, N11410);
nor NOR4 (N11421, N11415, N2937, N8095, N4484);
buf BUF1 (N11422, N11412);
buf BUF1 (N11423, N11421);
buf BUF1 (N11424, N11413);
buf BUF1 (N11425, N11423);
nand NAND4 (N11426, N11418, N10071, N2570, N8202);
not NOT1 (N11427, N11382);
xor XOR2 (N11428, N11420, N10399);
and AND3 (N11429, N11417, N679, N10962);
xor XOR2 (N11430, N11428, N510);
not NOT1 (N11431, N11427);
nand NAND3 (N11432, N11414, N8446, N7457);
buf BUF1 (N11433, N11432);
nand NAND4 (N11434, N11433, N8428, N7497, N3619);
not NOT1 (N11435, N11434);
or OR3 (N11436, N11426, N5091, N5093);
nor NOR2 (N11437, N11435, N1075);
or OR2 (N11438, N11419, N8403);
and AND3 (N11439, N11429, N9269, N10153);
nor NOR4 (N11440, N11439, N10503, N10438, N2630);
nor NOR2 (N11441, N11431, N9912);
nor NOR3 (N11442, N11438, N961, N2711);
or OR4 (N11443, N11403, N7273, N6949, N6534);
nor NOR4 (N11444, N11425, N116, N4767, N1742);
or OR3 (N11445, N11442, N3573, N1728);
and AND3 (N11446, N11437, N3240, N3378);
buf BUF1 (N11447, N11445);
xor XOR2 (N11448, N11446, N7368);
and AND2 (N11449, N11430, N6802);
and AND2 (N11450, N11424, N10915);
or OR2 (N11451, N11448, N6383);
not NOT1 (N11452, N11444);
nand NAND3 (N11453, N11436, N11164, N4251);
not NOT1 (N11454, N11449);
xor XOR2 (N11455, N11454, N1832);
or OR3 (N11456, N11452, N228, N467);
xor XOR2 (N11457, N11447, N4308);
buf BUF1 (N11458, N11456);
and AND3 (N11459, N11453, N6144, N253);
or OR3 (N11460, N11455, N6263, N1984);
or OR3 (N11461, N11458, N2249, N6684);
buf BUF1 (N11462, N11440);
and AND2 (N11463, N11443, N7860);
nor NOR4 (N11464, N11457, N1559, N8885, N2081);
nand NAND2 (N11465, N11422, N9935);
not NOT1 (N11466, N11459);
buf BUF1 (N11467, N11466);
xor XOR2 (N11468, N11464, N10610);
not NOT1 (N11469, N11441);
nand NAND2 (N11470, N11462, N1897);
nor NOR4 (N11471, N11463, N11244, N395, N4536);
or OR2 (N11472, N11471, N3734);
not NOT1 (N11473, N11460);
nand NAND4 (N11474, N11469, N9503, N515, N5446);
buf BUF1 (N11475, N11451);
nor NOR4 (N11476, N11472, N1915, N2609, N7330);
or OR3 (N11477, N11476, N6892, N10749);
not NOT1 (N11478, N11477);
and AND2 (N11479, N11475, N1131);
nor NOR3 (N11480, N11478, N11398, N9948);
buf BUF1 (N11481, N11480);
xor XOR2 (N11482, N11473, N8951);
and AND2 (N11483, N11461, N11422);
nor NOR2 (N11484, N11479, N8082);
xor XOR2 (N11485, N11465, N10838);
not NOT1 (N11486, N11468);
nor NOR3 (N11487, N11481, N1327, N8325);
nor NOR2 (N11488, N11484, N2975);
nor NOR3 (N11489, N11486, N2558, N11351);
nor NOR3 (N11490, N11487, N2646, N4468);
xor XOR2 (N11491, N11482, N7357);
or OR4 (N11492, N11490, N6154, N1800, N11031);
buf BUF1 (N11493, N11450);
nor NOR3 (N11494, N11493, N2653, N934);
or OR3 (N11495, N11491, N3257, N1158);
nor NOR4 (N11496, N11494, N7171, N5897, N6752);
or OR4 (N11497, N11485, N9200, N2483, N8507);
buf BUF1 (N11498, N11496);
buf BUF1 (N11499, N11492);
and AND2 (N11500, N11499, N3796);
or OR2 (N11501, N11497, N5787);
nand NAND4 (N11502, N11495, N1821, N11243, N8716);
xor XOR2 (N11503, N11500, N3278);
not NOT1 (N11504, N11489);
and AND2 (N11505, N11501, N6998);
nand NAND3 (N11506, N11488, N193, N3722);
nand NAND3 (N11507, N11474, N7084, N1079);
xor XOR2 (N11508, N11467, N3591);
or OR2 (N11509, N11508, N7687);
and AND4 (N11510, N11506, N6759, N584, N3416);
not NOT1 (N11511, N11498);
not NOT1 (N11512, N11510);
buf BUF1 (N11513, N11470);
nand NAND3 (N11514, N11503, N7091, N1899);
and AND3 (N11515, N11502, N3706, N8194);
and AND2 (N11516, N11514, N6157);
and AND3 (N11517, N11504, N6121, N9000);
not NOT1 (N11518, N11516);
nand NAND4 (N11519, N11507, N3977, N3102, N1094);
buf BUF1 (N11520, N11509);
not NOT1 (N11521, N11520);
and AND2 (N11522, N11517, N8524);
not NOT1 (N11523, N11483);
nor NOR4 (N11524, N11522, N624, N2175, N11257);
and AND3 (N11525, N11513, N2067, N6981);
or OR3 (N11526, N11525, N6569, N6607);
and AND2 (N11527, N11521, N424);
xor XOR2 (N11528, N11511, N5838);
nand NAND2 (N11529, N11518, N4459);
or OR2 (N11530, N11523, N4227);
xor XOR2 (N11531, N11519, N5121);
buf BUF1 (N11532, N11531);
xor XOR2 (N11533, N11524, N2240);
or OR4 (N11534, N11512, N776, N676, N6107);
xor XOR2 (N11535, N11530, N5097);
nor NOR3 (N11536, N11533, N9924, N8503);
nand NAND4 (N11537, N11534, N134, N10719, N1472);
xor XOR2 (N11538, N11532, N9136);
or OR3 (N11539, N11536, N10062, N6127);
xor XOR2 (N11540, N11539, N8220);
buf BUF1 (N11541, N11538);
xor XOR2 (N11542, N11526, N6937);
nor NOR4 (N11543, N11541, N9336, N6224, N2848);
and AND3 (N11544, N11529, N9400, N4702);
buf BUF1 (N11545, N11535);
buf BUF1 (N11546, N11543);
nand NAND4 (N11547, N11505, N5099, N2355, N5630);
not NOT1 (N11548, N11527);
nand NAND4 (N11549, N11547, N5990, N9583, N9831);
buf BUF1 (N11550, N11545);
and AND2 (N11551, N11515, N10854);
nand NAND4 (N11552, N11551, N3947, N2391, N361);
and AND2 (N11553, N11528, N1002);
or OR4 (N11554, N11548, N5585, N8562, N1283);
not NOT1 (N11555, N11553);
or OR4 (N11556, N11537, N2805, N9435, N789);
and AND2 (N11557, N11555, N8137);
nand NAND3 (N11558, N11542, N8572, N7854);
buf BUF1 (N11559, N11552);
nand NAND2 (N11560, N11558, N6215);
and AND2 (N11561, N11557, N6586);
nand NAND3 (N11562, N11540, N8964, N1713);
nand NAND3 (N11563, N11561, N5387, N9714);
and AND3 (N11564, N11562, N7105, N11276);
xor XOR2 (N11565, N11546, N2304);
xor XOR2 (N11566, N11549, N1020);
nor NOR2 (N11567, N11563, N6502);
nor NOR2 (N11568, N11565, N3858);
xor XOR2 (N11569, N11554, N10027);
not NOT1 (N11570, N11560);
nor NOR2 (N11571, N11570, N647);
nor NOR2 (N11572, N11567, N657);
not NOT1 (N11573, N11569);
and AND2 (N11574, N11572, N999);
and AND3 (N11575, N11550, N4482, N10434);
nand NAND4 (N11576, N11559, N985, N10219, N8620);
nor NOR2 (N11577, N11556, N11528);
not NOT1 (N11578, N11544);
nand NAND3 (N11579, N11575, N3998, N7704);
nor NOR2 (N11580, N11566, N11202);
buf BUF1 (N11581, N11568);
nand NAND4 (N11582, N11581, N7817, N6943, N10202);
or OR2 (N11583, N11580, N4369);
or OR2 (N11584, N11574, N11425);
nand NAND2 (N11585, N11582, N10923);
nor NOR3 (N11586, N11573, N3282, N8533);
buf BUF1 (N11587, N11583);
not NOT1 (N11588, N11564);
buf BUF1 (N11589, N11585);
nor NOR4 (N11590, N11578, N1448, N1560, N4485);
or OR2 (N11591, N11571, N3214);
and AND3 (N11592, N11586, N4410, N4455);
nor NOR3 (N11593, N11589, N1478, N1907);
buf BUF1 (N11594, N11587);
or OR4 (N11595, N11592, N2335, N3125, N7336);
nor NOR4 (N11596, N11591, N2129, N8329, N673);
buf BUF1 (N11597, N11576);
xor XOR2 (N11598, N11577, N2649);
or OR3 (N11599, N11588, N5541, N8861);
nor NOR3 (N11600, N11597, N206, N6588);
not NOT1 (N11601, N11590);
nand NAND2 (N11602, N11594, N9660);
or OR2 (N11603, N11595, N11414);
buf BUF1 (N11604, N11584);
nor NOR4 (N11605, N11596, N5945, N3336, N5021);
nor NOR3 (N11606, N11598, N6073, N1244);
buf BUF1 (N11607, N11602);
or OR2 (N11608, N11604, N1876);
or OR2 (N11609, N11605, N9021);
not NOT1 (N11610, N11606);
nand NAND4 (N11611, N11601, N10507, N11384, N5492);
buf BUF1 (N11612, N11600);
buf BUF1 (N11613, N11579);
buf BUF1 (N11614, N11612);
nand NAND4 (N11615, N11609, N6757, N7882, N2445);
buf BUF1 (N11616, N11614);
and AND4 (N11617, N11608, N3728, N3370, N9269);
nand NAND3 (N11618, N11603, N4414, N4428);
or OR3 (N11619, N11611, N1871, N2700);
nor NOR3 (N11620, N11619, N5976, N783);
not NOT1 (N11621, N11613);
or OR2 (N11622, N11593, N9862);
or OR4 (N11623, N11607, N2474, N2990, N8661);
nand NAND2 (N11624, N11618, N8162);
not NOT1 (N11625, N11624);
xor XOR2 (N11626, N11625, N2099);
and AND4 (N11627, N11621, N8854, N10955, N414);
nand NAND4 (N11628, N11620, N2444, N1562, N10278);
buf BUF1 (N11629, N11615);
not NOT1 (N11630, N11622);
nor NOR4 (N11631, N11599, N8125, N1428, N7280);
not NOT1 (N11632, N11616);
nand NAND3 (N11633, N11626, N4917, N3852);
or OR3 (N11634, N11628, N7062, N5888);
or OR2 (N11635, N11623, N9691);
nand NAND3 (N11636, N11617, N6767, N11236);
xor XOR2 (N11637, N11630, N7173);
or OR3 (N11638, N11610, N9146, N5365);
nand NAND2 (N11639, N11629, N1636);
buf BUF1 (N11640, N11631);
buf BUF1 (N11641, N11635);
xor XOR2 (N11642, N11634, N5842);
nor NOR2 (N11643, N11637, N5933);
nor NOR2 (N11644, N11639, N6214);
xor XOR2 (N11645, N11627, N9919);
buf BUF1 (N11646, N11640);
nand NAND2 (N11647, N11645, N7634);
nand NAND3 (N11648, N11632, N2730, N3171);
and AND4 (N11649, N11646, N218, N2842, N701);
xor XOR2 (N11650, N11638, N7389);
or OR3 (N11651, N11641, N3904, N8496);
or OR3 (N11652, N11633, N3344, N986);
and AND4 (N11653, N11648, N2053, N6723, N8428);
nand NAND4 (N11654, N11650, N6924, N7128, N7236);
xor XOR2 (N11655, N11653, N5203);
buf BUF1 (N11656, N11654);
nand NAND3 (N11657, N11656, N7705, N8458);
buf BUF1 (N11658, N11647);
nor NOR3 (N11659, N11651, N8372, N11632);
nor NOR3 (N11660, N11659, N6750, N7127);
and AND4 (N11661, N11652, N2540, N1271, N1573);
and AND4 (N11662, N11636, N2262, N11642, N1441);
not NOT1 (N11663, N7530);
not NOT1 (N11664, N11655);
buf BUF1 (N11665, N11661);
and AND4 (N11666, N11664, N7790, N4152, N6532);
nand NAND3 (N11667, N11649, N9869, N6366);
not NOT1 (N11668, N11658);
or OR2 (N11669, N11660, N265);
xor XOR2 (N11670, N11657, N718);
and AND4 (N11671, N11643, N11143, N1660, N9847);
nor NOR4 (N11672, N11663, N857, N3287, N9296);
nand NAND2 (N11673, N11669, N2321);
or OR4 (N11674, N11662, N6774, N4384, N3545);
and AND3 (N11675, N11671, N7613, N3696);
and AND2 (N11676, N11666, N6442);
xor XOR2 (N11677, N11665, N5569);
nand NAND2 (N11678, N11676, N7741);
buf BUF1 (N11679, N11673);
xor XOR2 (N11680, N11678, N1592);
or OR4 (N11681, N11667, N9532, N4583, N9587);
or OR2 (N11682, N11668, N1800);
nand NAND3 (N11683, N11675, N10667, N10133);
nor NOR4 (N11684, N11681, N4781, N9658, N2185);
nand NAND4 (N11685, N11683, N4560, N7138, N2979);
and AND3 (N11686, N11679, N2199, N10929);
buf BUF1 (N11687, N11680);
or OR3 (N11688, N11672, N9731, N10386);
nand NAND4 (N11689, N11686, N11615, N825, N315);
nor NOR3 (N11690, N11674, N1888, N9259);
nand NAND4 (N11691, N11687, N2750, N6079, N10798);
not NOT1 (N11692, N11684);
and AND4 (N11693, N11685, N2443, N3425, N2113);
buf BUF1 (N11694, N11693);
buf BUF1 (N11695, N11670);
xor XOR2 (N11696, N11677, N308);
xor XOR2 (N11697, N11690, N9528);
nor NOR4 (N11698, N11644, N5771, N4837, N6001);
buf BUF1 (N11699, N11689);
or OR4 (N11700, N11694, N3740, N3299, N302);
buf BUF1 (N11701, N11682);
and AND4 (N11702, N11695, N3137, N7121, N7464);
not NOT1 (N11703, N11688);
nand NAND2 (N11704, N11696, N2934);
or OR2 (N11705, N11704, N9649);
or OR3 (N11706, N11701, N5346, N4921);
buf BUF1 (N11707, N11692);
buf BUF1 (N11708, N11703);
and AND2 (N11709, N11697, N8922);
or OR2 (N11710, N11691, N2484);
buf BUF1 (N11711, N11709);
xor XOR2 (N11712, N11708, N6893);
xor XOR2 (N11713, N11707, N9918);
nand NAND4 (N11714, N11711, N9009, N2268, N5618);
xor XOR2 (N11715, N11698, N5109);
not NOT1 (N11716, N11715);
not NOT1 (N11717, N11713);
not NOT1 (N11718, N11705);
or OR4 (N11719, N11716, N11537, N6589, N3454);
nor NOR3 (N11720, N11719, N6854, N5932);
nand NAND3 (N11721, N11706, N11554, N9634);
nor NOR3 (N11722, N11717, N3592, N2700);
nand NAND2 (N11723, N11718, N9097);
xor XOR2 (N11724, N11723, N11167);
nor NOR2 (N11725, N11724, N2457);
nand NAND2 (N11726, N11700, N185);
buf BUF1 (N11727, N11712);
buf BUF1 (N11728, N11726);
or OR3 (N11729, N11725, N3842, N8603);
not NOT1 (N11730, N11729);
nor NOR3 (N11731, N11730, N643, N4);
nor NOR3 (N11732, N11720, N8765, N10660);
or OR3 (N11733, N11722, N5737, N9344);
not NOT1 (N11734, N11699);
nor NOR4 (N11735, N11728, N6601, N4097, N4694);
not NOT1 (N11736, N11734);
nor NOR2 (N11737, N11714, N9276);
nand NAND3 (N11738, N11733, N10140, N4680);
nor NOR2 (N11739, N11731, N1725);
nor NOR3 (N11740, N11737, N4501, N8590);
or OR3 (N11741, N11739, N4204, N5814);
and AND2 (N11742, N11736, N6688);
xor XOR2 (N11743, N11741, N10784);
not NOT1 (N11744, N11740);
nand NAND3 (N11745, N11710, N4650, N6506);
nor NOR3 (N11746, N11732, N902, N5995);
or OR3 (N11747, N11721, N11262, N632);
not NOT1 (N11748, N11747);
or OR3 (N11749, N11735, N2894, N3163);
not NOT1 (N11750, N11743);
xor XOR2 (N11751, N11702, N3409);
nand NAND4 (N11752, N11749, N513, N9107, N4026);
not NOT1 (N11753, N11748);
nor NOR2 (N11754, N11753, N7858);
buf BUF1 (N11755, N11750);
and AND4 (N11756, N11751, N6644, N11505, N6650);
xor XOR2 (N11757, N11756, N2029);
buf BUF1 (N11758, N11738);
not NOT1 (N11759, N11754);
xor XOR2 (N11760, N11744, N5512);
or OR3 (N11761, N11760, N2285, N1948);
or OR4 (N11762, N11759, N10755, N11258, N10209);
not NOT1 (N11763, N11757);
not NOT1 (N11764, N11758);
xor XOR2 (N11765, N11755, N6737);
and AND3 (N11766, N11765, N10656, N746);
buf BUF1 (N11767, N11752);
or OR4 (N11768, N11746, N8874, N4415, N9494);
and AND3 (N11769, N11767, N6019, N6957);
nor NOR3 (N11770, N11745, N5911, N1792);
not NOT1 (N11771, N11766);
nor NOR2 (N11772, N11762, N6589);
nor NOR3 (N11773, N11771, N7878, N1934);
not NOT1 (N11774, N11772);
nor NOR4 (N11775, N11727, N4494, N11724, N4987);
and AND3 (N11776, N11742, N8770, N8178);
not NOT1 (N11777, N11774);
xor XOR2 (N11778, N11764, N7298);
nand NAND2 (N11779, N11773, N1938);
nor NOR4 (N11780, N11779, N8780, N8668, N11433);
not NOT1 (N11781, N11777);
and AND2 (N11782, N11768, N7833);
xor XOR2 (N11783, N11776, N10092);
xor XOR2 (N11784, N11783, N10163);
nor NOR4 (N11785, N11763, N4705, N11675, N552);
xor XOR2 (N11786, N11775, N8461);
buf BUF1 (N11787, N11782);
nor NOR4 (N11788, N11770, N4175, N7670, N5313);
or OR2 (N11789, N11785, N10328);
or OR3 (N11790, N11761, N2790, N2753);
buf BUF1 (N11791, N11780);
not NOT1 (N11792, N11789);
or OR2 (N11793, N11787, N9443);
not NOT1 (N11794, N11791);
nor NOR3 (N11795, N11778, N2357, N8724);
or OR2 (N11796, N11781, N11244);
nand NAND4 (N11797, N11784, N4564, N1009, N6225);
buf BUF1 (N11798, N11769);
nor NOR4 (N11799, N11795, N6998, N5395, N7168);
nor NOR3 (N11800, N11792, N7722, N11065);
or OR4 (N11801, N11786, N6887, N6346, N11250);
not NOT1 (N11802, N11788);
nand NAND2 (N11803, N11802, N2755);
or OR2 (N11804, N11794, N4252);
nand NAND3 (N11805, N11804, N9125, N4591);
xor XOR2 (N11806, N11800, N3769);
xor XOR2 (N11807, N11803, N8491);
or OR2 (N11808, N11799, N8405);
and AND4 (N11809, N11793, N6081, N3436, N8707);
nor NOR3 (N11810, N11801, N10005, N2527);
not NOT1 (N11811, N11805);
nor NOR3 (N11812, N11809, N9989, N8230);
not NOT1 (N11813, N11811);
buf BUF1 (N11814, N11810);
or OR2 (N11815, N11798, N7011);
buf BUF1 (N11816, N11796);
or OR4 (N11817, N11807, N1201, N2611, N1415);
or OR2 (N11818, N11808, N7034);
buf BUF1 (N11819, N11818);
and AND3 (N11820, N11816, N2844, N147);
buf BUF1 (N11821, N11815);
nand NAND3 (N11822, N11806, N10872, N1203);
and AND2 (N11823, N11817, N10411);
or OR2 (N11824, N11797, N278);
or OR4 (N11825, N11823, N3183, N11664, N166);
not NOT1 (N11826, N11790);
or OR4 (N11827, N11814, N7784, N729, N6140);
xor XOR2 (N11828, N11822, N1903);
or OR4 (N11829, N11826, N6319, N10446, N8453);
nand NAND2 (N11830, N11812, N4217);
nor NOR2 (N11831, N11825, N8296);
or OR4 (N11832, N11820, N1242, N9543, N11096);
not NOT1 (N11833, N11819);
buf BUF1 (N11834, N11833);
nand NAND3 (N11835, N11821, N6709, N3159);
not NOT1 (N11836, N11824);
and AND2 (N11837, N11832, N2592);
not NOT1 (N11838, N11831);
or OR2 (N11839, N11837, N700);
nor NOR2 (N11840, N11838, N8469);
nand NAND3 (N11841, N11829, N8104, N6379);
not NOT1 (N11842, N11830);
nor NOR4 (N11843, N11840, N8127, N4839, N1611);
nor NOR3 (N11844, N11839, N2629, N3137);
and AND2 (N11845, N11828, N4296);
and AND4 (N11846, N11843, N10586, N3861, N1450);
nor NOR3 (N11847, N11835, N1454, N4908);
or OR3 (N11848, N11813, N11273, N7917);
xor XOR2 (N11849, N11848, N5841);
not NOT1 (N11850, N11844);
xor XOR2 (N11851, N11846, N4552);
nor NOR2 (N11852, N11834, N9108);
nand NAND3 (N11853, N11851, N7535, N6191);
and AND3 (N11854, N11845, N11156, N1536);
buf BUF1 (N11855, N11849);
or OR3 (N11856, N11827, N11687, N8547);
or OR2 (N11857, N11856, N4880);
buf BUF1 (N11858, N11850);
buf BUF1 (N11859, N11836);
xor XOR2 (N11860, N11841, N3045);
xor XOR2 (N11861, N11858, N6371);
and AND3 (N11862, N11861, N5498, N2296);
nand NAND2 (N11863, N11852, N291);
not NOT1 (N11864, N11854);
or OR4 (N11865, N11855, N2724, N2330, N5332);
and AND4 (N11866, N11847, N3829, N8496, N10067);
buf BUF1 (N11867, N11842);
nor NOR3 (N11868, N11857, N741, N10984);
and AND4 (N11869, N11866, N7183, N8790, N5461);
or OR3 (N11870, N11860, N5612, N4755);
or OR3 (N11871, N11862, N10364, N1901);
and AND2 (N11872, N11863, N6095);
xor XOR2 (N11873, N11868, N1576);
or OR3 (N11874, N11870, N6442, N4901);
buf BUF1 (N11875, N11864);
xor XOR2 (N11876, N11875, N6580);
nand NAND4 (N11877, N11873, N6467, N5718, N6176);
nor NOR3 (N11878, N11865, N11013, N4458);
buf BUF1 (N11879, N11853);
not NOT1 (N11880, N11879);
or OR4 (N11881, N11874, N6744, N6260, N11105);
xor XOR2 (N11882, N11878, N425);
or OR3 (N11883, N11880, N4648, N2488);
or OR4 (N11884, N11881, N4097, N4751, N10094);
and AND2 (N11885, N11876, N6091);
buf BUF1 (N11886, N11871);
nand NAND4 (N11887, N11886, N6478, N10170, N9828);
or OR4 (N11888, N11859, N3854, N6555, N6481);
not NOT1 (N11889, N11887);
or OR4 (N11890, N11885, N11549, N141, N1825);
buf BUF1 (N11891, N11888);
nor NOR3 (N11892, N11889, N7104, N10261);
nand NAND3 (N11893, N11884, N2988, N4532);
buf BUF1 (N11894, N11893);
not NOT1 (N11895, N11891);
buf BUF1 (N11896, N11882);
not NOT1 (N11897, N11896);
xor XOR2 (N11898, N11897, N3591);
nand NAND2 (N11899, N11890, N8242);
and AND2 (N11900, N11877, N2396);
not NOT1 (N11901, N11872);
nand NAND4 (N11902, N11899, N412, N6496, N8750);
or OR3 (N11903, N11895, N2116, N8103);
xor XOR2 (N11904, N11892, N3270);
or OR2 (N11905, N11894, N6692);
buf BUF1 (N11906, N11883);
nor NOR3 (N11907, N11900, N10341, N4207);
nand NAND3 (N11908, N11898, N3806, N11265);
or OR2 (N11909, N11901, N3896);
nand NAND4 (N11910, N11867, N7044, N3681, N55);
buf BUF1 (N11911, N11869);
nor NOR2 (N11912, N11909, N3358);
not NOT1 (N11913, N11904);
and AND4 (N11914, N11911, N206, N7945, N933);
buf BUF1 (N11915, N11908);
and AND2 (N11916, N11907, N5399);
buf BUF1 (N11917, N11910);
or OR3 (N11918, N11903, N11354, N3082);
nor NOR4 (N11919, N11914, N8763, N9886, N706);
and AND3 (N11920, N11918, N10276, N1170);
buf BUF1 (N11921, N11920);
xor XOR2 (N11922, N11919, N5712);
buf BUF1 (N11923, N11921);
or OR3 (N11924, N11922, N3747, N1195);
xor XOR2 (N11925, N11924, N10878);
xor XOR2 (N11926, N11923, N10722);
xor XOR2 (N11927, N11916, N2823);
xor XOR2 (N11928, N11912, N4130);
xor XOR2 (N11929, N11928, N10991);
buf BUF1 (N11930, N11906);
nand NAND4 (N11931, N11915, N3568, N2613, N3771);
nand NAND4 (N11932, N11902, N11805, N5861, N272);
nand NAND3 (N11933, N11930, N3320, N4469);
and AND2 (N11934, N11932, N6772);
nor NOR4 (N11935, N11925, N8577, N4297, N5180);
and AND2 (N11936, N11933, N7720);
not NOT1 (N11937, N11935);
or OR2 (N11938, N11929, N9145);
not NOT1 (N11939, N11936);
nor NOR2 (N11940, N11938, N7386);
or OR3 (N11941, N11927, N559, N231);
not NOT1 (N11942, N11940);
or OR3 (N11943, N11939, N9388, N130);
nor NOR2 (N11944, N11943, N3002);
nand NAND3 (N11945, N11931, N2436, N8291);
and AND3 (N11946, N11934, N11164, N1670);
and AND4 (N11947, N11941, N3246, N121, N8323);
nand NAND3 (N11948, N11905, N6070, N2305);
or OR4 (N11949, N11937, N7520, N159, N5914);
nor NOR3 (N11950, N11945, N6583, N11191);
xor XOR2 (N11951, N11948, N8798);
buf BUF1 (N11952, N11942);
nand NAND4 (N11953, N11949, N2935, N6813, N10571);
nand NAND3 (N11954, N11946, N1903, N7077);
or OR2 (N11955, N11951, N697);
not NOT1 (N11956, N11954);
and AND3 (N11957, N11950, N5562, N7260);
nand NAND4 (N11958, N11955, N10838, N9716, N4255);
not NOT1 (N11959, N11957);
or OR3 (N11960, N11917, N853, N467);
buf BUF1 (N11961, N11960);
xor XOR2 (N11962, N11958, N7394);
nor NOR3 (N11963, N11961, N168, N1949);
not NOT1 (N11964, N11963);
or OR2 (N11965, N11953, N10887);
buf BUF1 (N11966, N11947);
nor NOR2 (N11967, N11913, N9605);
nand NAND4 (N11968, N11966, N3124, N1465, N9505);
buf BUF1 (N11969, N11962);
or OR3 (N11970, N11952, N8277, N8074);
not NOT1 (N11971, N11969);
or OR4 (N11972, N11926, N4185, N4667, N7281);
nor NOR4 (N11973, N11968, N2974, N5774, N10814);
or OR3 (N11974, N11972, N5900, N8585);
nor NOR3 (N11975, N11970, N9539, N7304);
not NOT1 (N11976, N11964);
and AND4 (N11977, N11971, N9877, N4431, N7006);
nand NAND4 (N11978, N11965, N3773, N5591, N11581);
not NOT1 (N11979, N11977);
xor XOR2 (N11980, N11976, N1001);
not NOT1 (N11981, N11980);
nor NOR3 (N11982, N11975, N2224, N2998);
buf BUF1 (N11983, N11979);
nor NOR3 (N11984, N11983, N11472, N7756);
buf BUF1 (N11985, N11981);
not NOT1 (N11986, N11956);
buf BUF1 (N11987, N11959);
and AND3 (N11988, N11986, N3135, N11497);
and AND2 (N11989, N11974, N2173);
nor NOR3 (N11990, N11985, N7354, N514);
nand NAND3 (N11991, N11988, N2880, N10697);
xor XOR2 (N11992, N11982, N9633);
nor NOR2 (N11993, N11992, N11136);
not NOT1 (N11994, N11973);
not NOT1 (N11995, N11967);
nand NAND3 (N11996, N11987, N291, N4126);
nand NAND3 (N11997, N11989, N11419, N7253);
buf BUF1 (N11998, N11996);
buf BUF1 (N11999, N11997);
buf BUF1 (N12000, N11994);
buf BUF1 (N12001, N11991);
nand NAND2 (N12002, N11990, N10589);
xor XOR2 (N12003, N11998, N4454);
nor NOR4 (N12004, N11999, N2130, N2545, N4488);
nor NOR4 (N12005, N11993, N5108, N11110, N5902);
and AND2 (N12006, N11995, N10460);
and AND3 (N12007, N12006, N1966, N5847);
nand NAND3 (N12008, N11984, N5302, N9087);
buf BUF1 (N12009, N12002);
and AND4 (N12010, N12004, N3240, N10695, N11642);
nor NOR3 (N12011, N12008, N1394, N2403);
and AND2 (N12012, N11978, N382);
nor NOR3 (N12013, N12009, N7434, N6969);
nor NOR2 (N12014, N12012, N8997);
nand NAND3 (N12015, N12005, N7001, N3588);
and AND2 (N12016, N12007, N3393);
not NOT1 (N12017, N12015);
nand NAND4 (N12018, N12014, N11059, N1020, N3265);
nor NOR3 (N12019, N12001, N2954, N4299);
nand NAND2 (N12020, N12017, N10071);
nor NOR2 (N12021, N12003, N5770);
xor XOR2 (N12022, N12011, N5122);
or OR2 (N12023, N12020, N7876);
and AND4 (N12024, N12018, N716, N11653, N7848);
and AND4 (N12025, N12021, N1568, N6715, N4645);
nor NOR2 (N12026, N12023, N11071);
xor XOR2 (N12027, N12024, N6866);
not NOT1 (N12028, N12010);
nor NOR3 (N12029, N12026, N5421, N9271);
and AND4 (N12030, N12019, N10716, N3218, N4883);
or OR3 (N12031, N12013, N4785, N754);
nor NOR2 (N12032, N12029, N1579);
or OR2 (N12033, N12030, N7644);
buf BUF1 (N12034, N12016);
nor NOR3 (N12035, N11944, N2925, N302);
xor XOR2 (N12036, N12027, N11193);
xor XOR2 (N12037, N12025, N6801);
and AND3 (N12038, N12036, N8273, N11753);
nor NOR2 (N12039, N12035, N1579);
nor NOR3 (N12040, N12034, N3010, N11704);
not NOT1 (N12041, N12038);
not NOT1 (N12042, N12039);
nor NOR2 (N12043, N12037, N9835);
buf BUF1 (N12044, N12033);
or OR4 (N12045, N12022, N8331, N10192, N11615);
xor XOR2 (N12046, N12028, N6565);
nor NOR2 (N12047, N12041, N7833);
buf BUF1 (N12048, N12045);
xor XOR2 (N12049, N12032, N11020);
and AND3 (N12050, N12046, N4975, N11704);
or OR3 (N12051, N12031, N4929, N8458);
nor NOR4 (N12052, N12049, N10007, N7916, N7049);
and AND3 (N12053, N12050, N1694, N3885);
not NOT1 (N12054, N12052);
buf BUF1 (N12055, N12047);
xor XOR2 (N12056, N12054, N11125);
or OR4 (N12057, N12000, N10438, N11523, N9795);
nor NOR4 (N12058, N12044, N4924, N2039, N10036);
nand NAND3 (N12059, N12053, N7529, N5702);
or OR4 (N12060, N12057, N944, N4615, N7568);
or OR3 (N12061, N12051, N5169, N1719);
nand NAND4 (N12062, N12061, N10095, N867, N756);
nor NOR4 (N12063, N12060, N1643, N6836, N8153);
buf BUF1 (N12064, N12040);
not NOT1 (N12065, N12055);
xor XOR2 (N12066, N12043, N2257);
or OR2 (N12067, N12058, N6359);
nand NAND4 (N12068, N12059, N1255, N7341, N2435);
nor NOR2 (N12069, N12065, N4698);
nor NOR4 (N12070, N12069, N10591, N11187, N8805);
buf BUF1 (N12071, N12056);
nor NOR4 (N12072, N12063, N6315, N8958, N6059);
nand NAND4 (N12073, N12072, N4907, N6545, N8811);
buf BUF1 (N12074, N12073);
or OR4 (N12075, N12062, N9637, N8830, N346);
buf BUF1 (N12076, N12074);
buf BUF1 (N12077, N12070);
buf BUF1 (N12078, N12048);
nand NAND3 (N12079, N12071, N11689, N8059);
buf BUF1 (N12080, N12079);
or OR2 (N12081, N12080, N506);
xor XOR2 (N12082, N12077, N4274);
xor XOR2 (N12083, N12066, N12040);
and AND2 (N12084, N12042, N10894);
and AND4 (N12085, N12068, N6931, N3162, N10476);
nand NAND2 (N12086, N12082, N1781);
nand NAND4 (N12087, N12067, N11804, N10966, N1300);
nand NAND3 (N12088, N12085, N7941, N7132);
nand NAND2 (N12089, N12087, N7793);
nand NAND3 (N12090, N12089, N7058, N2401);
and AND2 (N12091, N12078, N4043);
not NOT1 (N12092, N12064);
nor NOR4 (N12093, N12084, N11266, N3732, N9478);
or OR2 (N12094, N12086, N5491);
or OR4 (N12095, N12076, N10820, N2190, N7628);
nor NOR4 (N12096, N12095, N3819, N4598, N4500);
and AND2 (N12097, N12096, N2405);
buf BUF1 (N12098, N12075);
and AND3 (N12099, N12093, N5204, N1221);
or OR4 (N12100, N12091, N3109, N3136, N11105);
not NOT1 (N12101, N12097);
or OR2 (N12102, N12100, N3475);
nand NAND3 (N12103, N12092, N956, N4926);
nand NAND3 (N12104, N12083, N7763, N2706);
nor NOR2 (N12105, N12099, N2812);
nand NAND2 (N12106, N12101, N7735);
buf BUF1 (N12107, N12104);
buf BUF1 (N12108, N12090);
nand NAND3 (N12109, N12105, N6601, N9738);
nor NOR2 (N12110, N12109, N6238);
nor NOR4 (N12111, N12102, N10836, N7159, N11597);
not NOT1 (N12112, N12108);
nor NOR4 (N12113, N12081, N7436, N10568, N8539);
and AND2 (N12114, N12107, N6350);
and AND4 (N12115, N12114, N8302, N8250, N9099);
or OR4 (N12116, N12103, N9816, N10143, N10339);
nand NAND2 (N12117, N12112, N7607);
or OR2 (N12118, N12094, N3758);
xor XOR2 (N12119, N12115, N2144);
xor XOR2 (N12120, N12110, N858);
xor XOR2 (N12121, N12119, N8881);
xor XOR2 (N12122, N12117, N1765);
buf BUF1 (N12123, N12111);
not NOT1 (N12124, N12118);
not NOT1 (N12125, N12124);
nor NOR2 (N12126, N12122, N2567);
buf BUF1 (N12127, N12125);
and AND2 (N12128, N12123, N5482);
nand NAND3 (N12129, N12121, N1173, N753);
xor XOR2 (N12130, N12126, N7367);
nor NOR3 (N12131, N12098, N57, N74);
and AND2 (N12132, N12113, N7298);
xor XOR2 (N12133, N12131, N5885);
buf BUF1 (N12134, N12120);
nor NOR4 (N12135, N12127, N8821, N3970, N5864);
and AND2 (N12136, N12128, N6860);
nor NOR2 (N12137, N12116, N1338);
nand NAND2 (N12138, N12136, N4979);
or OR2 (N12139, N12134, N2120);
nor NOR3 (N12140, N12106, N10425, N2143);
xor XOR2 (N12141, N12129, N10390);
nand NAND2 (N12142, N12140, N1393);
buf BUF1 (N12143, N12130);
nand NAND2 (N12144, N12142, N11918);
not NOT1 (N12145, N12132);
not NOT1 (N12146, N12145);
nor NOR4 (N12147, N12137, N1815, N11221, N6952);
xor XOR2 (N12148, N12143, N6104);
nand NAND4 (N12149, N12139, N8807, N6821, N9051);
nand NAND4 (N12150, N12146, N7332, N11830, N481);
not NOT1 (N12151, N12135);
nand NAND3 (N12152, N12133, N57, N12084);
not NOT1 (N12153, N12151);
nand NAND3 (N12154, N12148, N10418, N4081);
not NOT1 (N12155, N12152);
or OR2 (N12156, N12155, N11316);
xor XOR2 (N12157, N12154, N10741);
or OR4 (N12158, N12088, N4615, N2820, N4665);
and AND4 (N12159, N12149, N11362, N7726, N11973);
xor XOR2 (N12160, N12150, N9583);
xor XOR2 (N12161, N12158, N3963);
and AND3 (N12162, N12156, N9099, N411);
nand NAND2 (N12163, N12153, N1288);
not NOT1 (N12164, N12162);
not NOT1 (N12165, N12163);
xor XOR2 (N12166, N12159, N9043);
xor XOR2 (N12167, N12160, N5060);
xor XOR2 (N12168, N12166, N3862);
nor NOR4 (N12169, N12157, N9016, N2799, N5070);
nor NOR2 (N12170, N12169, N86);
not NOT1 (N12171, N12141);
or OR4 (N12172, N12167, N973, N11781, N1710);
buf BUF1 (N12173, N12172);
and AND3 (N12174, N12165, N2696, N10275);
nand NAND3 (N12175, N12171, N11796, N4495);
nor NOR4 (N12176, N12170, N11343, N1243, N7029);
or OR4 (N12177, N12164, N550, N11129, N11532);
not NOT1 (N12178, N12175);
buf BUF1 (N12179, N12147);
xor XOR2 (N12180, N12179, N4072);
not NOT1 (N12181, N12180);
nor NOR3 (N12182, N12174, N6542, N11226);
not NOT1 (N12183, N12182);
nor NOR2 (N12184, N12161, N11530);
or OR2 (N12185, N12184, N10000);
nor NOR2 (N12186, N12183, N7752);
not NOT1 (N12187, N12173);
nand NAND2 (N12188, N12181, N4518);
nor NOR4 (N12189, N12185, N1082, N11871, N8914);
not NOT1 (N12190, N12187);
buf BUF1 (N12191, N12176);
or OR3 (N12192, N12144, N1485, N5189);
nand NAND2 (N12193, N12191, N10949);
not NOT1 (N12194, N12186);
buf BUF1 (N12195, N12188);
xor XOR2 (N12196, N12177, N6905);
buf BUF1 (N12197, N12189);
xor XOR2 (N12198, N12190, N4264);
or OR4 (N12199, N12195, N11227, N8662, N8672);
or OR4 (N12200, N12198, N963, N12061, N576);
not NOT1 (N12201, N12200);
xor XOR2 (N12202, N12178, N10393);
or OR2 (N12203, N12197, N3);
nand NAND2 (N12204, N12168, N399);
not NOT1 (N12205, N12203);
nor NOR3 (N12206, N12201, N2924, N10152);
and AND4 (N12207, N12202, N2284, N4597, N10464);
and AND2 (N12208, N12206, N11786);
nor NOR4 (N12209, N12199, N7529, N6850, N5847);
nor NOR2 (N12210, N12196, N6598);
buf BUF1 (N12211, N12209);
buf BUF1 (N12212, N12208);
and AND3 (N12213, N12212, N4435, N4838);
not NOT1 (N12214, N12211);
and AND2 (N12215, N12214, N1553);
xor XOR2 (N12216, N12205, N2982);
or OR3 (N12217, N12210, N1205, N4907);
nand NAND2 (N12218, N12138, N5986);
nor NOR2 (N12219, N12213, N12022);
not NOT1 (N12220, N12207);
not NOT1 (N12221, N12192);
nor NOR2 (N12222, N12219, N8930);
not NOT1 (N12223, N12216);
or OR3 (N12224, N12194, N12031, N5415);
or OR2 (N12225, N12193, N4225);
nand NAND3 (N12226, N12220, N11625, N5044);
nand NAND3 (N12227, N12217, N6150, N2492);
buf BUF1 (N12228, N12221);
nor NOR2 (N12229, N12204, N10527);
nand NAND4 (N12230, N12229, N1140, N8478, N11889);
not NOT1 (N12231, N12227);
and AND2 (N12232, N12218, N5520);
xor XOR2 (N12233, N12230, N10441);
or OR2 (N12234, N12231, N9906);
nor NOR2 (N12235, N12226, N1701);
and AND4 (N12236, N12235, N10127, N7943, N1954);
nor NOR2 (N12237, N12232, N3266);
xor XOR2 (N12238, N12236, N1303);
not NOT1 (N12239, N12224);
xor XOR2 (N12240, N12238, N1522);
xor XOR2 (N12241, N12222, N10604);
nor NOR2 (N12242, N12234, N609);
and AND2 (N12243, N12233, N5098);
nand NAND3 (N12244, N12228, N11033, N12208);
buf BUF1 (N12245, N12237);
xor XOR2 (N12246, N12225, N2951);
buf BUF1 (N12247, N12245);
buf BUF1 (N12248, N12244);
nor NOR2 (N12249, N12223, N2492);
and AND4 (N12250, N12247, N3442, N2806, N657);
buf BUF1 (N12251, N12239);
nor NOR2 (N12252, N12241, N9665);
nor NOR4 (N12253, N12242, N9994, N9006, N3608);
nand NAND4 (N12254, N12240, N5966, N11227, N5356);
or OR4 (N12255, N12254, N6848, N1676, N9922);
nor NOR3 (N12256, N12246, N8285, N11439);
xor XOR2 (N12257, N12255, N3198);
and AND3 (N12258, N12257, N6664, N1386);
or OR4 (N12259, N12256, N4542, N11101, N10426);
buf BUF1 (N12260, N12253);
and AND4 (N12261, N12258, N6099, N8940, N1220);
nor NOR4 (N12262, N12252, N6311, N6613, N981);
and AND3 (N12263, N12243, N8653, N10974);
buf BUF1 (N12264, N12249);
buf BUF1 (N12265, N12264);
not NOT1 (N12266, N12260);
nand NAND4 (N12267, N12261, N1111, N4166, N4035);
nor NOR3 (N12268, N12266, N8039, N8530);
nand NAND2 (N12269, N12251, N4975);
not NOT1 (N12270, N12215);
buf BUF1 (N12271, N12259);
or OR3 (N12272, N12270, N86, N2305);
nor NOR2 (N12273, N12262, N11360);
buf BUF1 (N12274, N12248);
and AND2 (N12275, N12268, N2848);
and AND4 (N12276, N12269, N76, N8885, N6267);
and AND3 (N12277, N12267, N5930, N8527);
and AND3 (N12278, N12263, N10999, N2192);
and AND4 (N12279, N12276, N8170, N7127, N11126);
xor XOR2 (N12280, N12250, N3718);
or OR4 (N12281, N12277, N5500, N5437, N9835);
nor NOR4 (N12282, N12274, N3718, N487, N7068);
xor XOR2 (N12283, N12278, N10287);
nand NAND3 (N12284, N12283, N9688, N1732);
and AND3 (N12285, N12265, N4613, N7201);
xor XOR2 (N12286, N12279, N7848);
and AND3 (N12287, N12284, N10817, N3436);
buf BUF1 (N12288, N12273);
xor XOR2 (N12289, N12275, N5720);
and AND4 (N12290, N12288, N10281, N4251, N10909);
buf BUF1 (N12291, N12289);
buf BUF1 (N12292, N12285);
or OR2 (N12293, N12292, N11831);
nor NOR4 (N12294, N12281, N8252, N3985, N5147);
buf BUF1 (N12295, N12291);
and AND3 (N12296, N12282, N11344, N1074);
nor NOR4 (N12297, N12286, N7652, N8985, N9309);
or OR2 (N12298, N12296, N11845);
or OR4 (N12299, N12287, N9591, N2808, N7122);
xor XOR2 (N12300, N12294, N2883);
not NOT1 (N12301, N12297);
nand NAND3 (N12302, N12298, N5771, N3133);
xor XOR2 (N12303, N12272, N8933);
not NOT1 (N12304, N12271);
not NOT1 (N12305, N12299);
nor NOR2 (N12306, N12303, N7978);
nor NOR2 (N12307, N12295, N3723);
and AND2 (N12308, N12306, N11018);
and AND4 (N12309, N12302, N1087, N2060, N7648);
xor XOR2 (N12310, N12290, N5880);
buf BUF1 (N12311, N12309);
buf BUF1 (N12312, N12311);
nor NOR2 (N12313, N12293, N1170);
xor XOR2 (N12314, N12307, N3588);
buf BUF1 (N12315, N12305);
not NOT1 (N12316, N12310);
not NOT1 (N12317, N12300);
xor XOR2 (N12318, N12313, N5176);
nor NOR2 (N12319, N12280, N1138);
xor XOR2 (N12320, N12315, N6960);
not NOT1 (N12321, N12314);
xor XOR2 (N12322, N12318, N5272);
or OR4 (N12323, N12316, N2199, N4997, N940);
or OR4 (N12324, N12319, N10450, N7492, N5912);
buf BUF1 (N12325, N12323);
not NOT1 (N12326, N12322);
nand NAND4 (N12327, N12312, N4834, N3219, N7691);
not NOT1 (N12328, N12327);
and AND3 (N12329, N12328, N11423, N11896);
xor XOR2 (N12330, N12301, N1829);
nor NOR3 (N12331, N12321, N3411, N9248);
buf BUF1 (N12332, N12308);
or OR3 (N12333, N12332, N6085, N10037);
nor NOR4 (N12334, N12320, N2636, N9132, N6535);
not NOT1 (N12335, N12331);
nand NAND2 (N12336, N12330, N4773);
nand NAND4 (N12337, N12324, N8200, N8750, N5808);
buf BUF1 (N12338, N12329);
nor NOR3 (N12339, N12326, N4517, N2688);
nor NOR2 (N12340, N12317, N1840);
or OR2 (N12341, N12340, N3219);
or OR4 (N12342, N12341, N7351, N709, N10892);
buf BUF1 (N12343, N12333);
nor NOR3 (N12344, N12338, N6611, N6249);
or OR4 (N12345, N12325, N11848, N4958, N9986);
and AND3 (N12346, N12337, N6906, N3792);
or OR4 (N12347, N12346, N12044, N1359, N1434);
nand NAND3 (N12348, N12304, N8252, N1241);
and AND3 (N12349, N12336, N7709, N1129);
not NOT1 (N12350, N12334);
and AND3 (N12351, N12343, N2060, N1314);
not NOT1 (N12352, N12342);
xor XOR2 (N12353, N12344, N9538);
or OR4 (N12354, N12339, N7989, N6491, N5582);
or OR3 (N12355, N12347, N1899, N11986);
or OR3 (N12356, N12335, N5637, N11307);
or OR3 (N12357, N12352, N11901, N1066);
or OR4 (N12358, N12353, N11091, N3321, N11149);
nor NOR3 (N12359, N12355, N12326, N3502);
or OR3 (N12360, N12350, N4253, N9273);
xor XOR2 (N12361, N12357, N8934);
buf BUF1 (N12362, N12361);
nand NAND2 (N12363, N12348, N8450);
or OR3 (N12364, N12345, N11290, N10873);
xor XOR2 (N12365, N12354, N9464);
nor NOR3 (N12366, N12360, N6059, N12251);
not NOT1 (N12367, N12366);
buf BUF1 (N12368, N12364);
and AND4 (N12369, N12359, N11662, N2672, N12307);
buf BUF1 (N12370, N12356);
and AND3 (N12371, N12365, N8421, N7767);
or OR2 (N12372, N12370, N10162);
nor NOR4 (N12373, N12358, N2065, N1106, N5559);
buf BUF1 (N12374, N12368);
or OR2 (N12375, N12374, N3449);
xor XOR2 (N12376, N12351, N1181);
xor XOR2 (N12377, N12363, N11381);
xor XOR2 (N12378, N12375, N965);
xor XOR2 (N12379, N12362, N2671);
nor NOR3 (N12380, N12372, N11724, N7130);
and AND2 (N12381, N12373, N11139);
not NOT1 (N12382, N12377);
not NOT1 (N12383, N12369);
not NOT1 (N12384, N12378);
not NOT1 (N12385, N12382);
nand NAND2 (N12386, N12381, N2235);
nor NOR3 (N12387, N12386, N2786, N8838);
buf BUF1 (N12388, N12349);
buf BUF1 (N12389, N12379);
xor XOR2 (N12390, N12388, N2475);
or OR4 (N12391, N12367, N8087, N2662, N6290);
not NOT1 (N12392, N12376);
nand NAND3 (N12393, N12391, N2283, N5774);
not NOT1 (N12394, N12380);
not NOT1 (N12395, N12390);
buf BUF1 (N12396, N12385);
buf BUF1 (N12397, N12371);
or OR2 (N12398, N12387, N9552);
nor NOR2 (N12399, N12398, N764);
not NOT1 (N12400, N12393);
or OR4 (N12401, N12383, N9045, N3220, N11251);
nor NOR2 (N12402, N12394, N10918);
xor XOR2 (N12403, N12400, N9951);
nand NAND2 (N12404, N12396, N8635);
xor XOR2 (N12405, N12399, N11969);
and AND4 (N12406, N12397, N1679, N6846, N5873);
and AND3 (N12407, N12404, N4513, N8240);
nor NOR2 (N12408, N12405, N1968);
or OR4 (N12409, N12403, N11582, N7964, N10503);
xor XOR2 (N12410, N12409, N3277);
nand NAND4 (N12411, N12401, N2467, N7032, N1097);
buf BUF1 (N12412, N12407);
or OR3 (N12413, N12406, N7175, N4318);
nand NAND3 (N12414, N12412, N994, N10300);
not NOT1 (N12415, N12392);
xor XOR2 (N12416, N12402, N3185);
buf BUF1 (N12417, N12410);
xor XOR2 (N12418, N12395, N4629);
nor NOR2 (N12419, N12416, N5834);
nand NAND2 (N12420, N12389, N10951);
nor NOR3 (N12421, N12414, N12258, N11314);
buf BUF1 (N12422, N12419);
and AND3 (N12423, N12384, N6802, N5325);
buf BUF1 (N12424, N12408);
nand NAND4 (N12425, N12418, N2081, N6166, N3774);
nor NOR4 (N12426, N12421, N618, N10196, N125);
and AND2 (N12427, N12426, N6527);
nor NOR2 (N12428, N12425, N3378);
nand NAND2 (N12429, N12423, N12035);
nand NAND3 (N12430, N12427, N8498, N11934);
nor NOR4 (N12431, N12417, N10581, N6382, N2077);
buf BUF1 (N12432, N12415);
xor XOR2 (N12433, N12430, N9910);
nor NOR4 (N12434, N12420, N678, N1443, N2824);
nor NOR4 (N12435, N12433, N10464, N5104, N9500);
not NOT1 (N12436, N12422);
not NOT1 (N12437, N12435);
nor NOR2 (N12438, N12428, N8534);
nor NOR3 (N12439, N12429, N4554, N2502);
or OR4 (N12440, N12431, N4984, N569, N12041);
nand NAND3 (N12441, N12432, N2415, N10062);
buf BUF1 (N12442, N12441);
nor NOR2 (N12443, N12442, N9834);
and AND4 (N12444, N12443, N11890, N10004, N797);
nor NOR3 (N12445, N12438, N314, N3588);
nor NOR3 (N12446, N12445, N2943, N3759);
nor NOR3 (N12447, N12424, N6803, N7148);
buf BUF1 (N12448, N12413);
not NOT1 (N12449, N12411);
buf BUF1 (N12450, N12437);
xor XOR2 (N12451, N12439, N4222);
xor XOR2 (N12452, N12449, N6291);
buf BUF1 (N12453, N12434);
nand NAND3 (N12454, N12446, N4801, N8378);
xor XOR2 (N12455, N12451, N9564);
not NOT1 (N12456, N12440);
and AND4 (N12457, N12453, N7028, N10664, N7590);
nand NAND2 (N12458, N12454, N11908);
nor NOR2 (N12459, N12450, N11628);
and AND2 (N12460, N12458, N7050);
xor XOR2 (N12461, N12459, N10289);
not NOT1 (N12462, N12460);
nand NAND4 (N12463, N12462, N6361, N5664, N4825);
and AND4 (N12464, N12463, N3224, N8913, N9378);
nor NOR2 (N12465, N12452, N4908);
and AND2 (N12466, N12444, N8649);
and AND3 (N12467, N12456, N5597, N5225);
nor NOR3 (N12468, N12467, N4383, N11597);
not NOT1 (N12469, N12448);
and AND3 (N12470, N12447, N9006, N12262);
and AND3 (N12471, N12461, N10277, N11471);
not NOT1 (N12472, N12457);
nor NOR4 (N12473, N12470, N2897, N4054, N11760);
xor XOR2 (N12474, N12455, N5306);
and AND3 (N12475, N12474, N5581, N3820);
or OR3 (N12476, N12472, N1892, N211);
nor NOR2 (N12477, N12475, N11030);
xor XOR2 (N12478, N12477, N4820);
buf BUF1 (N12479, N12468);
nor NOR2 (N12480, N12479, N9732);
not NOT1 (N12481, N12473);
xor XOR2 (N12482, N12478, N6841);
or OR2 (N12483, N12481, N9407);
nand NAND2 (N12484, N12466, N8758);
and AND2 (N12485, N12482, N5338);
nor NOR4 (N12486, N12436, N160, N7091, N9800);
xor XOR2 (N12487, N12483, N628);
xor XOR2 (N12488, N12465, N5845);
or OR4 (N12489, N12484, N6356, N6266, N12052);
xor XOR2 (N12490, N12485, N4477);
nor NOR3 (N12491, N12469, N5646, N3960);
buf BUF1 (N12492, N12471);
nand NAND2 (N12493, N12480, N3063);
not NOT1 (N12494, N12490);
nand NAND3 (N12495, N12491, N2249, N3693);
nand NAND2 (N12496, N12488, N388);
nand NAND3 (N12497, N12489, N7095, N1783);
nand NAND2 (N12498, N12494, N10645);
nand NAND4 (N12499, N12492, N3689, N1173, N9562);
not NOT1 (N12500, N12487);
nor NOR3 (N12501, N12476, N11831, N3206);
or OR4 (N12502, N12496, N2608, N10506, N3873);
and AND4 (N12503, N12497, N5756, N11557, N3313);
nor NOR3 (N12504, N12464, N10700, N7523);
or OR3 (N12505, N12499, N8508, N4053);
not NOT1 (N12506, N12504);
or OR2 (N12507, N12493, N9883);
xor XOR2 (N12508, N12486, N7796);
and AND3 (N12509, N12495, N6490, N11253);
nand NAND3 (N12510, N12503, N12276, N3654);
nor NOR2 (N12511, N12502, N444);
not NOT1 (N12512, N12507);
xor XOR2 (N12513, N12506, N4750);
buf BUF1 (N12514, N12498);
nor NOR3 (N12515, N12505, N902, N8564);
xor XOR2 (N12516, N12501, N6152);
or OR2 (N12517, N12515, N229);
buf BUF1 (N12518, N12510);
or OR3 (N12519, N12516, N6261, N9788);
nor NOR3 (N12520, N12517, N8437, N4902);
or OR2 (N12521, N12520, N10206);
nor NOR2 (N12522, N12500, N8763);
nor NOR3 (N12523, N12511, N5157, N8196);
and AND3 (N12524, N12514, N7047, N931);
not NOT1 (N12525, N12512);
buf BUF1 (N12526, N12521);
and AND2 (N12527, N12519, N428);
buf BUF1 (N12528, N12518);
not NOT1 (N12529, N12524);
nor NOR3 (N12530, N12513, N4040, N8575);
or OR2 (N12531, N12523, N1867);
and AND2 (N12532, N12530, N12346);
buf BUF1 (N12533, N12508);
and AND4 (N12534, N12509, N6768, N7810, N9783);
xor XOR2 (N12535, N12527, N4520);
and AND2 (N12536, N12534, N10068);
and AND4 (N12537, N12525, N3138, N2481, N870);
xor XOR2 (N12538, N12532, N2966);
nand NAND3 (N12539, N12529, N2666, N8753);
buf BUF1 (N12540, N12535);
and AND4 (N12541, N12537, N1519, N4649, N11350);
xor XOR2 (N12542, N12538, N10011);
buf BUF1 (N12543, N12526);
nor NOR2 (N12544, N12540, N3043);
and AND2 (N12545, N12544, N9292);
nand NAND3 (N12546, N12541, N3911, N12425);
buf BUF1 (N12547, N12543);
and AND4 (N12548, N12545, N4696, N8368, N5819);
not NOT1 (N12549, N12528);
nand NAND4 (N12550, N12533, N4253, N6280, N12414);
not NOT1 (N12551, N12522);
nand NAND4 (N12552, N12550, N297, N10327, N777);
nand NAND3 (N12553, N12531, N4888, N10359);
nor NOR4 (N12554, N12539, N10475, N9620, N4421);
and AND4 (N12555, N12551, N694, N9591, N12521);
or OR4 (N12556, N12547, N2840, N9978, N8326);
nor NOR3 (N12557, N12555, N8310, N2038);
nor NOR4 (N12558, N12552, N7274, N9966, N513);
or OR4 (N12559, N12553, N11961, N2745, N11985);
buf BUF1 (N12560, N12549);
nor NOR3 (N12561, N12556, N267, N5495);
xor XOR2 (N12562, N12554, N7072);
xor XOR2 (N12563, N12562, N1845);
nand NAND4 (N12564, N12548, N1774, N6964, N10808);
or OR4 (N12565, N12557, N12092, N6621, N10204);
buf BUF1 (N12566, N12561);
nor NOR2 (N12567, N12546, N6553);
nand NAND3 (N12568, N12564, N10835, N11292);
xor XOR2 (N12569, N12565, N2180);
nand NAND3 (N12570, N12536, N2340, N1784);
buf BUF1 (N12571, N12559);
xor XOR2 (N12572, N12566, N85);
and AND3 (N12573, N12569, N2905, N5819);
and AND3 (N12574, N12558, N4093, N7204);
nand NAND3 (N12575, N12560, N2290, N2995);
and AND4 (N12576, N12542, N10667, N11813, N3868);
not NOT1 (N12577, N12576);
and AND4 (N12578, N12567, N5133, N9470, N9229);
xor XOR2 (N12579, N12577, N6333);
or OR3 (N12580, N12578, N2998, N1200);
nor NOR3 (N12581, N12575, N8187, N2390);
nor NOR2 (N12582, N12572, N8770);
and AND2 (N12583, N12582, N9436);
xor XOR2 (N12584, N12579, N8362);
nand NAND3 (N12585, N12584, N1659, N4950);
not NOT1 (N12586, N12571);
buf BUF1 (N12587, N12574);
nor NOR3 (N12588, N12587, N3907, N8809);
buf BUF1 (N12589, N12586);
nor NOR3 (N12590, N12568, N5159, N3114);
nand NAND3 (N12591, N12589, N7604, N5847);
nand NAND3 (N12592, N12591, N12169, N11623);
xor XOR2 (N12593, N12590, N7438);
not NOT1 (N12594, N12580);
nand NAND4 (N12595, N12583, N12138, N8096, N12489);
xor XOR2 (N12596, N12594, N3965);
buf BUF1 (N12597, N12595);
xor XOR2 (N12598, N12596, N12415);
nor NOR2 (N12599, N12563, N11899);
or OR2 (N12600, N12597, N5502);
not NOT1 (N12601, N12592);
nor NOR3 (N12602, N12593, N4504, N5347);
or OR4 (N12603, N12581, N7066, N10849, N4520);
nand NAND4 (N12604, N12602, N5792, N10228, N5420);
nor NOR3 (N12605, N12600, N11641, N10079);
nand NAND4 (N12606, N12570, N347, N7490, N7411);
and AND2 (N12607, N12601, N2049);
nor NOR4 (N12608, N12607, N11164, N7106, N8588);
nand NAND2 (N12609, N12608, N851);
nand NAND3 (N12610, N12599, N10289, N952);
and AND3 (N12611, N12603, N5768, N10401);
buf BUF1 (N12612, N12610);
buf BUF1 (N12613, N12604);
or OR3 (N12614, N12609, N3527, N8504);
nand NAND2 (N12615, N12613, N3436);
buf BUF1 (N12616, N12614);
or OR4 (N12617, N12598, N11048, N7073, N8560);
nor NOR4 (N12618, N12588, N6905, N8002, N8769);
nor NOR2 (N12619, N12616, N8467);
nand NAND3 (N12620, N12617, N11624, N3157);
not NOT1 (N12621, N12585);
buf BUF1 (N12622, N12606);
buf BUF1 (N12623, N12619);
not NOT1 (N12624, N12620);
xor XOR2 (N12625, N12605, N7105);
nand NAND3 (N12626, N12623, N2041, N7210);
xor XOR2 (N12627, N12624, N12314);
or OR4 (N12628, N12625, N3752, N8615, N426);
nor NOR3 (N12629, N12627, N11748, N10705);
and AND3 (N12630, N12626, N516, N8201);
not NOT1 (N12631, N12612);
xor XOR2 (N12632, N12573, N365);
nor NOR2 (N12633, N12628, N5423);
and AND3 (N12634, N12615, N1276, N1450);
and AND2 (N12635, N12621, N10900);
xor XOR2 (N12636, N12634, N6451);
nand NAND2 (N12637, N12631, N10051);
nand NAND4 (N12638, N12637, N10504, N12621, N9577);
or OR2 (N12639, N12635, N10186);
nor NOR2 (N12640, N12630, N6846);
and AND4 (N12641, N12636, N9084, N11914, N2314);
xor XOR2 (N12642, N12638, N10668);
xor XOR2 (N12643, N12618, N6683);
buf BUF1 (N12644, N12640);
xor XOR2 (N12645, N12643, N915);
or OR2 (N12646, N12639, N11681);
xor XOR2 (N12647, N12611, N12368);
and AND3 (N12648, N12646, N1924, N6838);
and AND3 (N12649, N12642, N1286, N11812);
not NOT1 (N12650, N12632);
xor XOR2 (N12651, N12649, N5082);
buf BUF1 (N12652, N12650);
nand NAND2 (N12653, N12647, N373);
or OR3 (N12654, N12629, N7909, N10019);
nor NOR4 (N12655, N12633, N10029, N140, N4020);
nand NAND3 (N12656, N12653, N11368, N12313);
nand NAND3 (N12657, N12654, N2468, N6744);
and AND4 (N12658, N12644, N3917, N7727, N12567);
and AND4 (N12659, N12657, N3105, N5783, N4919);
nor NOR2 (N12660, N12655, N951);
buf BUF1 (N12661, N12641);
xor XOR2 (N12662, N12661, N3745);
and AND2 (N12663, N12645, N6015);
xor XOR2 (N12664, N12658, N1010);
xor XOR2 (N12665, N12660, N2296);
xor XOR2 (N12666, N12656, N6040);
not NOT1 (N12667, N12662);
not NOT1 (N12668, N12666);
buf BUF1 (N12669, N12659);
not NOT1 (N12670, N12668);
xor XOR2 (N12671, N12667, N694);
and AND2 (N12672, N12665, N6024);
nand NAND4 (N12673, N12652, N6575, N1028, N1543);
buf BUF1 (N12674, N12663);
or OR4 (N12675, N12670, N2489, N4444, N9013);
nor NOR2 (N12676, N12651, N5843);
xor XOR2 (N12677, N12622, N4988);
not NOT1 (N12678, N12669);
or OR2 (N12679, N12677, N10038);
not NOT1 (N12680, N12674);
and AND2 (N12681, N12678, N819);
buf BUF1 (N12682, N12679);
and AND2 (N12683, N12672, N12217);
and AND2 (N12684, N12675, N4804);
buf BUF1 (N12685, N12680);
not NOT1 (N12686, N12676);
not NOT1 (N12687, N12682);
nand NAND4 (N12688, N12684, N3727, N11292, N1440);
nor NOR2 (N12689, N12664, N7423);
buf BUF1 (N12690, N12673);
nand NAND3 (N12691, N12683, N2564, N8613);
nand NAND4 (N12692, N12685, N10206, N1763, N7311);
nor NOR3 (N12693, N12688, N2634, N1481);
or OR2 (N12694, N12691, N2938);
buf BUF1 (N12695, N12693);
not NOT1 (N12696, N12671);
nor NOR3 (N12697, N12690, N555, N8611);
and AND3 (N12698, N12648, N12363, N8398);
or OR2 (N12699, N12696, N10202);
nor NOR3 (N12700, N12681, N9157, N6821);
buf BUF1 (N12701, N12700);
nand NAND3 (N12702, N12699, N6658, N10045);
nor NOR3 (N12703, N12687, N11942, N2600);
nor NOR3 (N12704, N12686, N9962, N3246);
buf BUF1 (N12705, N12702);
nor NOR4 (N12706, N12695, N498, N11898, N1637);
buf BUF1 (N12707, N12706);
or OR4 (N12708, N12697, N10717, N7765, N1830);
nand NAND3 (N12709, N12694, N4836, N4997);
and AND4 (N12710, N12692, N8303, N8464, N11235);
xor XOR2 (N12711, N12698, N9264);
xor XOR2 (N12712, N12703, N4305);
xor XOR2 (N12713, N12711, N2108);
buf BUF1 (N12714, N12704);
xor XOR2 (N12715, N12701, N3965);
buf BUF1 (N12716, N12715);
buf BUF1 (N12717, N12712);
xor XOR2 (N12718, N12710, N10503);
buf BUF1 (N12719, N12713);
nor NOR4 (N12720, N12717, N5557, N9754, N10016);
xor XOR2 (N12721, N12718, N3749);
or OR4 (N12722, N12714, N3366, N1398, N10088);
buf BUF1 (N12723, N12722);
and AND2 (N12724, N12708, N1494);
not NOT1 (N12725, N12719);
xor XOR2 (N12726, N12725, N7127);
nor NOR2 (N12727, N12707, N9937);
not NOT1 (N12728, N12721);
nor NOR3 (N12729, N12689, N10831, N4560);
or OR4 (N12730, N12728, N7103, N10432, N573);
xor XOR2 (N12731, N12716, N49);
buf BUF1 (N12732, N12731);
buf BUF1 (N12733, N12730);
not NOT1 (N12734, N12720);
xor XOR2 (N12735, N12727, N1365);
not NOT1 (N12736, N12724);
and AND3 (N12737, N12709, N1276, N11110);
xor XOR2 (N12738, N12737, N5408);
nor NOR3 (N12739, N12733, N12344, N5634);
buf BUF1 (N12740, N12726);
xor XOR2 (N12741, N12729, N7442);
nand NAND3 (N12742, N12739, N6617, N3858);
not NOT1 (N12743, N12742);
and AND2 (N12744, N12705, N7551);
or OR4 (N12745, N12743, N10131, N12030, N9656);
xor XOR2 (N12746, N12734, N9222);
xor XOR2 (N12747, N12735, N8173);
xor XOR2 (N12748, N12723, N5690);
xor XOR2 (N12749, N12744, N2657);
nor NOR3 (N12750, N12746, N4673, N6531);
and AND2 (N12751, N12740, N7209);
nor NOR3 (N12752, N12732, N9034, N5616);
and AND3 (N12753, N12748, N12053, N11697);
xor XOR2 (N12754, N12738, N781);
nor NOR2 (N12755, N12753, N1596);
buf BUF1 (N12756, N12750);
not NOT1 (N12757, N12745);
nand NAND3 (N12758, N12756, N7633, N10075);
nor NOR4 (N12759, N12736, N3969, N3530, N8262);
nor NOR4 (N12760, N12749, N7476, N4966, N3863);
nand NAND3 (N12761, N12757, N6426, N2189);
xor XOR2 (N12762, N12752, N4389);
and AND3 (N12763, N12741, N3813, N741);
xor XOR2 (N12764, N12762, N27);
nand NAND4 (N12765, N12751, N83, N6613, N11776);
nand NAND2 (N12766, N12763, N10628);
xor XOR2 (N12767, N12759, N5033);
nand NAND4 (N12768, N12767, N5664, N4147, N2315);
or OR3 (N12769, N12755, N6887, N11676);
xor XOR2 (N12770, N12760, N12329);
or OR2 (N12771, N12764, N292);
or OR3 (N12772, N12761, N8183, N4957);
xor XOR2 (N12773, N12770, N7620);
nor NOR4 (N12774, N12758, N4048, N9676, N4040);
nand NAND2 (N12775, N12766, N7632);
and AND4 (N12776, N12768, N12444, N11706, N12372);
nor NOR2 (N12777, N12754, N6299);
or OR4 (N12778, N12774, N12027, N6378, N757);
nand NAND2 (N12779, N12747, N1404);
or OR3 (N12780, N12771, N7950, N10983);
xor XOR2 (N12781, N12776, N1289);
and AND4 (N12782, N12772, N8838, N3649, N9993);
and AND2 (N12783, N12782, N978);
not NOT1 (N12784, N12773);
and AND3 (N12785, N12777, N9888, N4319);
nor NOR2 (N12786, N12780, N11989);
nand NAND3 (N12787, N12779, N2867, N1619);
buf BUF1 (N12788, N12778);
or OR2 (N12789, N12775, N7737);
and AND4 (N12790, N12785, N411, N7900, N2983);
not NOT1 (N12791, N12769);
not NOT1 (N12792, N12791);
and AND4 (N12793, N12790, N3321, N743, N4299);
nand NAND3 (N12794, N12786, N2010, N4734);
or OR2 (N12795, N12784, N4804);
nand NAND2 (N12796, N12788, N10884);
and AND2 (N12797, N12795, N2305);
or OR2 (N12798, N12765, N5546);
or OR4 (N12799, N12794, N2457, N12792, N9862);
xor XOR2 (N12800, N230, N7998);
nand NAND3 (N12801, N12789, N3757, N10853);
nand NAND2 (N12802, N12781, N5079);
or OR2 (N12803, N12796, N11070);
nand NAND3 (N12804, N12793, N3981, N1430);
not NOT1 (N12805, N12799);
nor NOR2 (N12806, N12805, N9797);
nor NOR4 (N12807, N12783, N2872, N6780, N8566);
xor XOR2 (N12808, N12802, N5778);
nor NOR2 (N12809, N12808, N1382);
or OR2 (N12810, N12807, N11668);
and AND2 (N12811, N12787, N3555);
buf BUF1 (N12812, N12800);
and AND3 (N12813, N12797, N11756, N9386);
not NOT1 (N12814, N12810);
or OR4 (N12815, N12812, N3909, N10524, N2885);
xor XOR2 (N12816, N12804, N5668);
buf BUF1 (N12817, N12816);
not NOT1 (N12818, N12815);
nand NAND4 (N12819, N12811, N9635, N6173, N12818);
xor XOR2 (N12820, N2240, N2669);
or OR3 (N12821, N12819, N2623, N5867);
and AND3 (N12822, N12801, N1811, N10352);
not NOT1 (N12823, N12803);
and AND3 (N12824, N12814, N959, N5598);
not NOT1 (N12825, N12822);
and AND3 (N12826, N12809, N2203, N398);
or OR3 (N12827, N12824, N7363, N4054);
buf BUF1 (N12828, N12823);
and AND2 (N12829, N12813, N10526);
xor XOR2 (N12830, N12821, N11813);
not NOT1 (N12831, N12830);
xor XOR2 (N12832, N12806, N10879);
or OR2 (N12833, N12828, N7146);
and AND2 (N12834, N12798, N3150);
and AND2 (N12835, N12820, N10410);
not NOT1 (N12836, N12825);
xor XOR2 (N12837, N12836, N4103);
or OR2 (N12838, N12832, N2249);
xor XOR2 (N12839, N12837, N3948);
not NOT1 (N12840, N12839);
and AND3 (N12841, N12826, N11457, N10821);
or OR2 (N12842, N12834, N9932);
nand NAND2 (N12843, N12833, N8558);
nand NAND2 (N12844, N12829, N1872);
buf BUF1 (N12845, N12844);
and AND2 (N12846, N12845, N9594);
nand NAND3 (N12847, N12827, N7405, N11962);
and AND3 (N12848, N12831, N5400, N788);
buf BUF1 (N12849, N12842);
nor NOR3 (N12850, N12840, N10106, N6841);
nand NAND3 (N12851, N12843, N11754, N4362);
buf BUF1 (N12852, N12847);
not NOT1 (N12853, N12849);
buf BUF1 (N12854, N12852);
or OR3 (N12855, N12846, N12596, N9247);
and AND2 (N12856, N12848, N7063);
and AND4 (N12857, N12838, N4796, N9855, N6477);
nand NAND2 (N12858, N12854, N10073);
and AND3 (N12859, N12850, N6749, N8238);
buf BUF1 (N12860, N12856);
buf BUF1 (N12861, N12859);
nor NOR4 (N12862, N12853, N2759, N4070, N3356);
and AND4 (N12863, N12860, N7483, N6886, N4168);
nor NOR4 (N12864, N12861, N6690, N4681, N5578);
nor NOR4 (N12865, N12851, N6870, N7968, N3574);
xor XOR2 (N12866, N12857, N5716);
xor XOR2 (N12867, N12862, N7929);
buf BUF1 (N12868, N12835);
or OR4 (N12869, N12863, N7483, N5793, N544);
or OR4 (N12870, N12841, N85, N8585, N11183);
nand NAND3 (N12871, N12869, N9494, N4949);
not NOT1 (N12872, N12858);
or OR4 (N12873, N12870, N12178, N9264, N12863);
and AND4 (N12874, N12871, N11172, N2904, N2310);
and AND4 (N12875, N12817, N11730, N3765, N10566);
not NOT1 (N12876, N12867);
buf BUF1 (N12877, N12868);
nand NAND3 (N12878, N12874, N9596, N5489);
or OR2 (N12879, N12864, N6809);
nor NOR2 (N12880, N12873, N364);
buf BUF1 (N12881, N12878);
nand NAND3 (N12882, N12876, N117, N943);
and AND3 (N12883, N12879, N2563, N8136);
not NOT1 (N12884, N12883);
nand NAND2 (N12885, N12855, N7664);
and AND3 (N12886, N12875, N4476, N7457);
not NOT1 (N12887, N12877);
nand NAND2 (N12888, N12872, N9362);
not NOT1 (N12889, N12886);
or OR3 (N12890, N12889, N8483, N11250);
nor NOR2 (N12891, N12882, N12017);
nand NAND4 (N12892, N12885, N7478, N7337, N6213);
nand NAND2 (N12893, N12890, N850);
buf BUF1 (N12894, N12884);
nor NOR2 (N12895, N12891, N10493);
not NOT1 (N12896, N12887);
or OR2 (N12897, N12880, N11413);
and AND4 (N12898, N12888, N12216, N12347, N7203);
not NOT1 (N12899, N12866);
nand NAND2 (N12900, N12898, N12713);
nand NAND3 (N12901, N12897, N5590, N3393);
and AND2 (N12902, N12896, N5880);
or OR3 (N12903, N12892, N11834, N5389);
and AND3 (N12904, N12900, N11653, N10516);
nand NAND2 (N12905, N12902, N1037);
or OR4 (N12906, N12903, N6367, N8596, N6410);
buf BUF1 (N12907, N12881);
or OR4 (N12908, N12895, N10384, N1375, N7808);
not NOT1 (N12909, N12899);
nor NOR4 (N12910, N12901, N4045, N12649, N12881);
or OR3 (N12911, N12909, N802, N10988);
nand NAND4 (N12912, N12904, N7093, N3572, N9417);
xor XOR2 (N12913, N12893, N1473);
and AND2 (N12914, N12910, N10527);
buf BUF1 (N12915, N12865);
not NOT1 (N12916, N12913);
or OR3 (N12917, N12912, N7465, N11572);
buf BUF1 (N12918, N12916);
buf BUF1 (N12919, N12894);
and AND2 (N12920, N12919, N3914);
nand NAND4 (N12921, N12914, N7654, N4001, N8731);
and AND4 (N12922, N12918, N11171, N12305, N4792);
nand NAND3 (N12923, N12921, N12211, N6820);
or OR2 (N12924, N12917, N4373);
not NOT1 (N12925, N12911);
buf BUF1 (N12926, N12925);
xor XOR2 (N12927, N12920, N7541);
buf BUF1 (N12928, N12906);
nand NAND3 (N12929, N12927, N11168, N4957);
buf BUF1 (N12930, N12923);
xor XOR2 (N12931, N12922, N240);
and AND3 (N12932, N12928, N6412, N1131);
xor XOR2 (N12933, N12930, N526);
and AND4 (N12934, N12907, N11553, N3569, N7454);
not NOT1 (N12935, N12908);
not NOT1 (N12936, N12935);
buf BUF1 (N12937, N12929);
not NOT1 (N12938, N12932);
nand NAND4 (N12939, N12933, N3253, N12459, N10529);
not NOT1 (N12940, N12924);
nand NAND4 (N12941, N12915, N893, N1064, N226);
or OR2 (N12942, N12939, N101);
buf BUF1 (N12943, N12937);
not NOT1 (N12944, N12938);
xor XOR2 (N12945, N12942, N4620);
nor NOR2 (N12946, N12931, N4543);
xor XOR2 (N12947, N12936, N2008);
nand NAND3 (N12948, N12946, N2206, N12377);
and AND2 (N12949, N12948, N4335);
nor NOR4 (N12950, N12940, N5275, N1677, N2627);
or OR2 (N12951, N12926, N10000);
not NOT1 (N12952, N12950);
nand NAND4 (N12953, N12934, N232, N1323, N12834);
xor XOR2 (N12954, N12944, N12806);
nand NAND3 (N12955, N12905, N1996, N10429);
nand NAND4 (N12956, N12947, N4672, N1657, N2385);
or OR3 (N12957, N12952, N6202, N4694);
xor XOR2 (N12958, N12953, N11946);
buf BUF1 (N12959, N12956);
xor XOR2 (N12960, N12957, N10173);
nand NAND4 (N12961, N12949, N1854, N3504, N8020);
and AND4 (N12962, N12954, N5864, N626, N12379);
buf BUF1 (N12963, N12955);
or OR2 (N12964, N12951, N2793);
and AND4 (N12965, N12963, N5187, N272, N12526);
buf BUF1 (N12966, N12945);
or OR4 (N12967, N12961, N10554, N10848, N3374);
nor NOR3 (N12968, N12941, N4015, N6341);
not NOT1 (N12969, N12964);
xor XOR2 (N12970, N12960, N543);
buf BUF1 (N12971, N12970);
or OR3 (N12972, N12969, N10234, N8453);
or OR4 (N12973, N12971, N7277, N10675, N11411);
nand NAND2 (N12974, N12973, N12699);
and AND4 (N12975, N12959, N4424, N1979, N8128);
buf BUF1 (N12976, N12965);
and AND4 (N12977, N12976, N9565, N1629, N5903);
xor XOR2 (N12978, N12974, N11500);
xor XOR2 (N12979, N12972, N12816);
nor NOR3 (N12980, N12978, N1206, N10042);
not NOT1 (N12981, N12958);
or OR2 (N12982, N12975, N12226);
or OR2 (N12983, N12966, N9410);
xor XOR2 (N12984, N12981, N7239);
not NOT1 (N12985, N12982);
not NOT1 (N12986, N12980);
buf BUF1 (N12987, N12979);
not NOT1 (N12988, N12962);
nand NAND3 (N12989, N12987, N8510, N8185);
buf BUF1 (N12990, N12984);
or OR2 (N12991, N12986, N12215);
buf BUF1 (N12992, N12968);
nand NAND3 (N12993, N12992, N1374, N1233);
nand NAND4 (N12994, N12943, N2072, N1323, N11331);
buf BUF1 (N12995, N12991);
nand NAND2 (N12996, N12989, N10083);
or OR4 (N12997, N12994, N10439, N11375, N9837);
buf BUF1 (N12998, N12996);
or OR3 (N12999, N12988, N3982, N5686);
not NOT1 (N13000, N12985);
not NOT1 (N13001, N12967);
buf BUF1 (N13002, N12995);
buf BUF1 (N13003, N12997);
nand NAND3 (N13004, N12998, N5136, N2589);
nand NAND3 (N13005, N13002, N10255, N7826);
nand NAND3 (N13006, N13003, N3463, N8787);
buf BUF1 (N13007, N13004);
buf BUF1 (N13008, N12977);
nor NOR2 (N13009, N13001, N11530);
xor XOR2 (N13010, N13008, N2917);
xor XOR2 (N13011, N12999, N3988);
or OR3 (N13012, N13009, N5752, N681);
or OR3 (N13013, N13005, N9371, N9337);
nor NOR2 (N13014, N13000, N3666);
xor XOR2 (N13015, N12993, N2774);
and AND4 (N13016, N13013, N10795, N6565, N6807);
buf BUF1 (N13017, N13015);
buf BUF1 (N13018, N13010);
not NOT1 (N13019, N13007);
nand NAND4 (N13020, N13018, N1999, N8697, N3860);
nand NAND3 (N13021, N13020, N6977, N1394);
not NOT1 (N13022, N13014);
xor XOR2 (N13023, N13021, N1913);
nand NAND3 (N13024, N13019, N1797, N7558);
or OR4 (N13025, N13024, N6405, N155, N12569);
buf BUF1 (N13026, N12990);
and AND4 (N13027, N13012, N1047, N11069, N10468);
not NOT1 (N13028, N13016);
nor NOR4 (N13029, N13017, N1879, N1755, N2370);
buf BUF1 (N13030, N12983);
or OR2 (N13031, N13026, N2469);
and AND4 (N13032, N13029, N5367, N699, N5736);
or OR2 (N13033, N13022, N229);
nor NOR3 (N13034, N13031, N8515, N12642);
and AND4 (N13035, N13025, N1955, N10650, N3166);
nor NOR2 (N13036, N13023, N3465);
not NOT1 (N13037, N13028);
or OR2 (N13038, N13011, N2434);
or OR3 (N13039, N13037, N6017, N2753);
nand NAND3 (N13040, N13032, N2817, N2267);
not NOT1 (N13041, N13027);
and AND2 (N13042, N13038, N8323);
xor XOR2 (N13043, N13036, N7165);
or OR3 (N13044, N13040, N12360, N8559);
or OR3 (N13045, N13039, N11071, N12972);
not NOT1 (N13046, N13006);
nand NAND2 (N13047, N13034, N5596);
xor XOR2 (N13048, N13041, N1881);
and AND2 (N13049, N13030, N12868);
buf BUF1 (N13050, N13044);
and AND3 (N13051, N13033, N9196, N11260);
not NOT1 (N13052, N13051);
xor XOR2 (N13053, N13047, N8789);
xor XOR2 (N13054, N13043, N11364);
nand NAND2 (N13055, N13048, N10891);
nand NAND2 (N13056, N13050, N4182);
nand NAND2 (N13057, N13035, N8370);
not NOT1 (N13058, N13055);
nor NOR2 (N13059, N13056, N9722);
and AND3 (N13060, N13059, N1999, N920);
xor XOR2 (N13061, N13053, N6276);
nand NAND4 (N13062, N13061, N6969, N2387, N5144);
not NOT1 (N13063, N13045);
nor NOR2 (N13064, N13049, N12474);
xor XOR2 (N13065, N13052, N9282);
and AND4 (N13066, N13060, N3784, N7293, N9785);
and AND4 (N13067, N13063, N7847, N6209, N36);
xor XOR2 (N13068, N13057, N559);
buf BUF1 (N13069, N13067);
and AND2 (N13070, N13058, N1383);
nand NAND3 (N13071, N13066, N3425, N10592);
buf BUF1 (N13072, N13042);
nand NAND2 (N13073, N13069, N9301);
and AND2 (N13074, N13054, N10740);
nand NAND2 (N13075, N13068, N6465);
xor XOR2 (N13076, N13075, N7806);
xor XOR2 (N13077, N13072, N6394);
nand NAND3 (N13078, N13073, N544, N4409);
nor NOR4 (N13079, N13071, N6193, N215, N10030);
and AND3 (N13080, N13070, N3420, N12069);
buf BUF1 (N13081, N13078);
and AND2 (N13082, N13079, N11702);
not NOT1 (N13083, N13081);
and AND3 (N13084, N13046, N9679, N6391);
not NOT1 (N13085, N13082);
and AND4 (N13086, N13077, N97, N9420, N6891);
xor XOR2 (N13087, N13062, N8387);
and AND4 (N13088, N13086, N12048, N4349, N6055);
not NOT1 (N13089, N13084);
xor XOR2 (N13090, N13083, N11875);
buf BUF1 (N13091, N13090);
nor NOR4 (N13092, N13088, N9246, N11121, N9849);
or OR2 (N13093, N13087, N9188);
or OR4 (N13094, N13092, N6414, N544, N6710);
or OR3 (N13095, N13091, N2961, N2437);
and AND3 (N13096, N13095, N5585, N10018);
xor XOR2 (N13097, N13089, N6802);
nor NOR2 (N13098, N13076, N3989);
or OR2 (N13099, N13097, N7194);
or OR2 (N13100, N13085, N10641);
not NOT1 (N13101, N13093);
and AND2 (N13102, N13094, N74);
nor NOR4 (N13103, N13101, N9901, N2629, N6493);
or OR2 (N13104, N13096, N2953);
and AND2 (N13105, N13102, N9928);
not NOT1 (N13106, N13105);
nor NOR3 (N13107, N13099, N4855, N10036);
and AND4 (N13108, N13100, N3, N4335, N6150);
buf BUF1 (N13109, N13098);
not NOT1 (N13110, N13064);
xor XOR2 (N13111, N13065, N7476);
and AND4 (N13112, N13108, N5359, N1805, N6898);
or OR2 (N13113, N13080, N4222);
nand NAND4 (N13114, N13113, N10549, N4947, N2001);
and AND4 (N13115, N13112, N7515, N1730, N7090);
and AND4 (N13116, N13109, N3702, N4421, N9478);
or OR3 (N13117, N13111, N7198, N5960);
xor XOR2 (N13118, N13103, N8323);
nor NOR4 (N13119, N13117, N12488, N7086, N9565);
nand NAND4 (N13120, N13114, N3206, N12504, N11699);
buf BUF1 (N13121, N13106);
xor XOR2 (N13122, N13116, N7102);
xor XOR2 (N13123, N13107, N6029);
or OR3 (N13124, N13121, N6641, N13114);
not NOT1 (N13125, N13104);
and AND4 (N13126, N13124, N11209, N9347, N9785);
nor NOR3 (N13127, N13115, N12915, N1180);
buf BUF1 (N13128, N13125);
nand NAND3 (N13129, N13074, N2156, N10864);
buf BUF1 (N13130, N13110);
nand NAND3 (N13131, N13119, N10627, N4147);
buf BUF1 (N13132, N13126);
and AND2 (N13133, N13127, N4820);
or OR4 (N13134, N13122, N7619, N6899, N8198);
not NOT1 (N13135, N13129);
nand NAND3 (N13136, N13120, N4066, N1840);
nand NAND3 (N13137, N13133, N7511, N12538);
not NOT1 (N13138, N13130);
xor XOR2 (N13139, N13118, N9496);
xor XOR2 (N13140, N13139, N7559);
xor XOR2 (N13141, N13135, N6555);
or OR4 (N13142, N13138, N3203, N11707, N4512);
or OR3 (N13143, N13128, N11182, N7809);
xor XOR2 (N13144, N13134, N2975);
xor XOR2 (N13145, N13142, N12635);
or OR2 (N13146, N13136, N7703);
nor NOR2 (N13147, N13132, N2447);
not NOT1 (N13148, N13123);
xor XOR2 (N13149, N13140, N10924);
not NOT1 (N13150, N13147);
or OR3 (N13151, N13148, N2776, N1364);
and AND3 (N13152, N13149, N10529, N2576);
nand NAND4 (N13153, N13141, N1305, N5140, N7914);
not NOT1 (N13154, N13151);
nand NAND3 (N13155, N13143, N1693, N4434);
xor XOR2 (N13156, N13152, N9393);
not NOT1 (N13157, N13146);
nand NAND2 (N13158, N13155, N5293);
or OR2 (N13159, N13153, N7014);
buf BUF1 (N13160, N13158);
nand NAND4 (N13161, N13159, N2311, N9128, N10876);
buf BUF1 (N13162, N13161);
nand NAND3 (N13163, N13145, N6889, N1330);
and AND2 (N13164, N13156, N7312);
not NOT1 (N13165, N13131);
or OR4 (N13166, N13157, N12990, N10155, N7487);
or OR4 (N13167, N13166, N8600, N911, N5748);
nor NOR4 (N13168, N13137, N3815, N347, N10750);
xor XOR2 (N13169, N13167, N1080);
and AND3 (N13170, N13144, N4005, N1882);
nor NOR4 (N13171, N13168, N3450, N2609, N12061);
xor XOR2 (N13172, N13163, N6984);
not NOT1 (N13173, N13172);
nor NOR4 (N13174, N13165, N10409, N9372, N10450);
nor NOR3 (N13175, N13170, N1401, N7575);
buf BUF1 (N13176, N13169);
not NOT1 (N13177, N13171);
xor XOR2 (N13178, N13173, N6634);
buf BUF1 (N13179, N13176);
nand NAND3 (N13180, N13150, N4273, N12624);
not NOT1 (N13181, N13175);
or OR3 (N13182, N13177, N10520, N11115);
nor NOR2 (N13183, N13174, N8148);
or OR4 (N13184, N13182, N7087, N7238, N3988);
nor NOR3 (N13185, N13181, N6213, N11577);
nand NAND4 (N13186, N13164, N1548, N12583, N748);
nand NAND4 (N13187, N13183, N7416, N3704, N11434);
buf BUF1 (N13188, N13160);
and AND4 (N13189, N13187, N13096, N7511, N3065);
buf BUF1 (N13190, N13188);
and AND3 (N13191, N13154, N12853, N7599);
and AND3 (N13192, N13180, N1266, N7509);
not NOT1 (N13193, N13178);
buf BUF1 (N13194, N13191);
xor XOR2 (N13195, N13162, N12719);
or OR2 (N13196, N13193, N1060);
not NOT1 (N13197, N13189);
xor XOR2 (N13198, N13192, N10498);
and AND2 (N13199, N13198, N3284);
not NOT1 (N13200, N13194);
and AND3 (N13201, N13186, N8519, N6372);
buf BUF1 (N13202, N13197);
and AND2 (N13203, N13179, N5010);
and AND2 (N13204, N13185, N5581);
not NOT1 (N13205, N13199);
and AND4 (N13206, N13204, N8106, N409, N7606);
and AND3 (N13207, N13201, N907, N9620);
not NOT1 (N13208, N13190);
nand NAND2 (N13209, N13205, N12096);
nor NOR3 (N13210, N13207, N2100, N1350);
nor NOR3 (N13211, N13200, N5914, N1031);
and AND3 (N13212, N13210, N389, N12971);
nand NAND3 (N13213, N13212, N13207, N2840);
not NOT1 (N13214, N13184);
nor NOR4 (N13215, N13203, N1192, N8642, N7540);
and AND3 (N13216, N13214, N4277, N7017);
nor NOR4 (N13217, N13206, N3093, N5531, N4282);
or OR3 (N13218, N13215, N7699, N10285);
not NOT1 (N13219, N13196);
nor NOR3 (N13220, N13209, N8935, N2284);
nor NOR3 (N13221, N13208, N3576, N12707);
not NOT1 (N13222, N13211);
buf BUF1 (N13223, N13216);
nand NAND2 (N13224, N13222, N2627);
nor NOR2 (N13225, N13213, N13025);
buf BUF1 (N13226, N13195);
not NOT1 (N13227, N13219);
and AND2 (N13228, N13227, N5950);
or OR4 (N13229, N13225, N6643, N10724, N3772);
not NOT1 (N13230, N13226);
or OR4 (N13231, N13224, N5049, N11819, N3609);
nand NAND3 (N13232, N13220, N11599, N2718);
not NOT1 (N13233, N13228);
nand NAND4 (N13234, N13218, N10827, N7651, N1715);
nor NOR2 (N13235, N13217, N5450);
not NOT1 (N13236, N13232);
and AND2 (N13237, N13202, N3);
nand NAND2 (N13238, N13230, N3952);
or OR2 (N13239, N13221, N5868);
xor XOR2 (N13240, N13237, N8968);
nor NOR3 (N13241, N13231, N10531, N6358);
xor XOR2 (N13242, N13229, N11265);
not NOT1 (N13243, N13239);
nor NOR3 (N13244, N13236, N10990, N11961);
nor NOR2 (N13245, N13223, N1939);
and AND2 (N13246, N13238, N4939);
and AND4 (N13247, N13234, N12900, N7813, N4240);
nand NAND2 (N13248, N13245, N3356);
or OR2 (N13249, N13248, N6731);
nand NAND2 (N13250, N13247, N3638);
nand NAND3 (N13251, N13233, N13180, N10458);
and AND4 (N13252, N13246, N7741, N9695, N7395);
and AND2 (N13253, N13250, N7230);
or OR2 (N13254, N13249, N3474);
xor XOR2 (N13255, N13242, N11785);
xor XOR2 (N13256, N13255, N2368);
xor XOR2 (N13257, N13252, N10504);
nand NAND2 (N13258, N13257, N3156);
xor XOR2 (N13259, N13241, N8029);
xor XOR2 (N13260, N13259, N9674);
or OR4 (N13261, N13260, N4169, N6210, N1180);
and AND3 (N13262, N13256, N3921, N9053);
and AND4 (N13263, N13251, N6367, N8238, N4118);
and AND4 (N13264, N13262, N9898, N6771, N9264);
xor XOR2 (N13265, N13244, N12731);
not NOT1 (N13266, N13235);
or OR2 (N13267, N13265, N10202);
not NOT1 (N13268, N13240);
and AND2 (N13269, N13267, N406);
and AND3 (N13270, N13243, N2400, N1586);
nand NAND3 (N13271, N13253, N1590, N10557);
nand NAND3 (N13272, N13268, N7603, N1265);
xor XOR2 (N13273, N13270, N5671);
buf BUF1 (N13274, N13264);
nand NAND4 (N13275, N13263, N5798, N10948, N5270);
xor XOR2 (N13276, N13258, N1128);
and AND2 (N13277, N13276, N9622);
buf BUF1 (N13278, N13277);
or OR2 (N13279, N13272, N6490);
buf BUF1 (N13280, N13269);
not NOT1 (N13281, N13271);
and AND3 (N13282, N13279, N4796, N4438);
nand NAND3 (N13283, N13273, N10978, N5204);
buf BUF1 (N13284, N13282);
or OR3 (N13285, N13278, N12973, N8619);
nor NOR3 (N13286, N13285, N5359, N7616);
not NOT1 (N13287, N13266);
not NOT1 (N13288, N13286);
not NOT1 (N13289, N13274);
and AND4 (N13290, N13289, N11423, N164, N4493);
xor XOR2 (N13291, N13284, N13041);
nor NOR2 (N13292, N13281, N10220);
or OR2 (N13293, N13275, N7358);
not NOT1 (N13294, N13254);
nand NAND2 (N13295, N13283, N10311);
nor NOR2 (N13296, N13280, N5198);
nor NOR4 (N13297, N13293, N11858, N950, N8375);
nand NAND2 (N13298, N13297, N13249);
or OR4 (N13299, N13287, N3668, N10235, N3500);
not NOT1 (N13300, N13299);
nand NAND4 (N13301, N13291, N9974, N10740, N9750);
nand NAND2 (N13302, N13296, N6329);
buf BUF1 (N13303, N13261);
buf BUF1 (N13304, N13295);
or OR2 (N13305, N13300, N7880);
not NOT1 (N13306, N13301);
xor XOR2 (N13307, N13288, N8919);
nand NAND3 (N13308, N13292, N12294, N1710);
and AND4 (N13309, N13306, N6508, N7140, N4462);
and AND4 (N13310, N13305, N11659, N10659, N10373);
or OR3 (N13311, N13303, N2055, N3814);
nor NOR3 (N13312, N13290, N92, N5922);
not NOT1 (N13313, N13294);
not NOT1 (N13314, N13304);
xor XOR2 (N13315, N13311, N9318);
buf BUF1 (N13316, N13310);
nor NOR2 (N13317, N13315, N9950);
nand NAND4 (N13318, N13313, N8206, N10457, N10682);
and AND4 (N13319, N13316, N6244, N12922, N5891);
buf BUF1 (N13320, N13312);
not NOT1 (N13321, N13318);
or OR2 (N13322, N13307, N12782);
nor NOR4 (N13323, N13322, N9749, N10853, N2218);
xor XOR2 (N13324, N13317, N6500);
buf BUF1 (N13325, N13323);
or OR3 (N13326, N13324, N3933, N1397);
and AND3 (N13327, N13309, N4420, N12111);
xor XOR2 (N13328, N13314, N4481);
nand NAND4 (N13329, N13321, N5281, N2685, N5304);
and AND3 (N13330, N13325, N5182, N10768);
xor XOR2 (N13331, N13328, N4172);
not NOT1 (N13332, N13308);
not NOT1 (N13333, N13327);
nor NOR2 (N13334, N13319, N3601);
and AND4 (N13335, N13329, N3727, N1611, N498);
or OR4 (N13336, N13298, N1131, N4999, N8882);
nand NAND3 (N13337, N13320, N8167, N10260);
not NOT1 (N13338, N13331);
not NOT1 (N13339, N13332);
nor NOR3 (N13340, N13334, N12672, N8220);
nand NAND2 (N13341, N13339, N10337);
not NOT1 (N13342, N13340);
not NOT1 (N13343, N13337);
or OR4 (N13344, N13341, N10771, N2485, N5476);
and AND4 (N13345, N13335, N9833, N7071, N6180);
buf BUF1 (N13346, N13344);
not NOT1 (N13347, N13342);
nor NOR2 (N13348, N13336, N11179);
nor NOR4 (N13349, N13346, N10417, N9326, N4360);
buf BUF1 (N13350, N13326);
or OR3 (N13351, N13347, N10796, N10426);
nand NAND4 (N13352, N13348, N3892, N5130, N11133);
and AND2 (N13353, N13352, N5292);
buf BUF1 (N13354, N13343);
or OR3 (N13355, N13345, N2782, N12594);
and AND2 (N13356, N13330, N9075);
buf BUF1 (N13357, N13349);
and AND3 (N13358, N13333, N3530, N9524);
nor NOR3 (N13359, N13350, N10203, N4073);
nand NAND3 (N13360, N13351, N7101, N9386);
xor XOR2 (N13361, N13357, N10299);
nand NAND2 (N13362, N13355, N1029);
nand NAND2 (N13363, N13360, N363);
not NOT1 (N13364, N13359);
buf BUF1 (N13365, N13354);
xor XOR2 (N13366, N13361, N5413);
xor XOR2 (N13367, N13362, N11899);
nor NOR4 (N13368, N13338, N4982, N3043, N6844);
buf BUF1 (N13369, N13302);
or OR4 (N13370, N13368, N10493, N12645, N10788);
and AND4 (N13371, N13369, N8819, N1145, N9683);
nand NAND3 (N13372, N13358, N9218, N4875);
xor XOR2 (N13373, N13353, N8978);
and AND4 (N13374, N13365, N787, N5656, N5968);
nor NOR2 (N13375, N13372, N1841);
xor XOR2 (N13376, N13364, N9241);
xor XOR2 (N13377, N13363, N6910);
or OR2 (N13378, N13377, N10217);
buf BUF1 (N13379, N13366);
and AND2 (N13380, N13371, N6744);
and AND3 (N13381, N13374, N5627, N9817);
nor NOR3 (N13382, N13379, N3773, N5755);
nand NAND3 (N13383, N13382, N8326, N7635);
not NOT1 (N13384, N13375);
not NOT1 (N13385, N13367);
or OR4 (N13386, N13376, N2194, N9723, N6529);
nor NOR3 (N13387, N13383, N8401, N4221);
and AND2 (N13388, N13380, N10482);
nor NOR3 (N13389, N13388, N171, N9551);
or OR3 (N13390, N13385, N10774, N10786);
buf BUF1 (N13391, N13356);
and AND4 (N13392, N13386, N510, N12611, N12969);
not NOT1 (N13393, N13373);
nor NOR3 (N13394, N13381, N4435, N7472);
nor NOR3 (N13395, N13391, N11239, N3471);
nand NAND2 (N13396, N13394, N12620);
buf BUF1 (N13397, N13393);
buf BUF1 (N13398, N13397);
and AND4 (N13399, N13396, N6315, N2642, N3383);
nand NAND2 (N13400, N13370, N6346);
xor XOR2 (N13401, N13378, N606);
nor NOR4 (N13402, N13384, N7823, N12468, N10729);
buf BUF1 (N13403, N13400);
xor XOR2 (N13404, N13402, N2788);
not NOT1 (N13405, N13389);
not NOT1 (N13406, N13387);
buf BUF1 (N13407, N13398);
not NOT1 (N13408, N13404);
or OR2 (N13409, N13407, N4458);
or OR3 (N13410, N13399, N12543, N7939);
and AND4 (N13411, N13392, N13359, N5171, N8384);
buf BUF1 (N13412, N13403);
not NOT1 (N13413, N13401);
buf BUF1 (N13414, N13390);
nand NAND2 (N13415, N13409, N9300);
not NOT1 (N13416, N13410);
nand NAND3 (N13417, N13395, N12276, N6839);
nand NAND3 (N13418, N13416, N11905, N2020);
or OR2 (N13419, N13405, N1672);
or OR4 (N13420, N13415, N7491, N12329, N5165);
or OR2 (N13421, N13418, N10094);
and AND4 (N13422, N13417, N5681, N10220, N7693);
and AND4 (N13423, N13414, N7246, N7814, N5623);
and AND2 (N13424, N13423, N11987);
and AND3 (N13425, N13424, N340, N1979);
xor XOR2 (N13426, N13419, N12072);
or OR4 (N13427, N13408, N3381, N8837, N13372);
nor NOR2 (N13428, N13413, N34);
nand NAND4 (N13429, N13412, N3827, N10379, N8139);
buf BUF1 (N13430, N13420);
nor NOR3 (N13431, N13427, N11664, N9554);
nor NOR3 (N13432, N13425, N5345, N8821);
nand NAND3 (N13433, N13426, N4315, N11821);
or OR2 (N13434, N13430, N6789);
buf BUF1 (N13435, N13421);
xor XOR2 (N13436, N13432, N10587);
and AND2 (N13437, N13433, N8232);
buf BUF1 (N13438, N13431);
buf BUF1 (N13439, N13406);
nand NAND3 (N13440, N13439, N4622, N4891);
nand NAND2 (N13441, N13435, N5795);
buf BUF1 (N13442, N13437);
nand NAND4 (N13443, N13434, N11660, N11602, N674);
nor NOR2 (N13444, N13428, N10465);
or OR3 (N13445, N13438, N485, N5492);
nor NOR2 (N13446, N13442, N5114);
buf BUF1 (N13447, N13411);
or OR2 (N13448, N13436, N8840);
nor NOR3 (N13449, N13444, N10145, N3745);
nand NAND3 (N13450, N13422, N2696, N8212);
nand NAND2 (N13451, N13449, N3804);
and AND4 (N13452, N13429, N6211, N5273, N9501);
and AND2 (N13453, N13446, N1873);
nor NOR4 (N13454, N13448, N11882, N9510, N7806);
buf BUF1 (N13455, N13454);
xor XOR2 (N13456, N13455, N12711);
nand NAND2 (N13457, N13451, N9391);
nor NOR2 (N13458, N13456, N4369);
buf BUF1 (N13459, N13440);
nand NAND3 (N13460, N13458, N10582, N1813);
or OR3 (N13461, N13459, N2048, N1764);
and AND3 (N13462, N13457, N11906, N2025);
not NOT1 (N13463, N13447);
nand NAND2 (N13464, N13441, N3895);
nand NAND3 (N13465, N13452, N7124, N746);
or OR3 (N13466, N13445, N13045, N4323);
not NOT1 (N13467, N13453);
and AND3 (N13468, N13467, N10203, N11062);
buf BUF1 (N13469, N13464);
nand NAND2 (N13470, N13466, N3229);
and AND3 (N13471, N13461, N3933, N10165);
or OR3 (N13472, N13463, N8534, N8400);
nand NAND3 (N13473, N13470, N11852, N11656);
or OR3 (N13474, N13450, N13288, N11582);
or OR4 (N13475, N13469, N78, N7247, N8208);
and AND4 (N13476, N13473, N5588, N7251, N12734);
nand NAND2 (N13477, N13476, N4910);
not NOT1 (N13478, N13468);
not NOT1 (N13479, N13443);
nor NOR3 (N13480, N13477, N11295, N9173);
buf BUF1 (N13481, N13471);
nor NOR4 (N13482, N13479, N3968, N2285, N10074);
nor NOR4 (N13483, N13480, N4809, N9871, N2579);
or OR2 (N13484, N13460, N8032);
nor NOR2 (N13485, N13481, N13278);
xor XOR2 (N13486, N13482, N7524);
nor NOR4 (N13487, N13472, N4397, N2281, N12933);
buf BUF1 (N13488, N13475);
xor XOR2 (N13489, N13488, N3986);
xor XOR2 (N13490, N13487, N9621);
xor XOR2 (N13491, N13483, N6055);
xor XOR2 (N13492, N13490, N11880);
or OR3 (N13493, N13489, N1096, N9886);
nor NOR3 (N13494, N13491, N11065, N3554);
or OR3 (N13495, N13494, N5781, N8071);
or OR4 (N13496, N13465, N10345, N1745, N2394);
and AND2 (N13497, N13484, N10064);
not NOT1 (N13498, N13485);
and AND2 (N13499, N13462, N4807);
nor NOR2 (N13500, N13499, N3071);
or OR4 (N13501, N13497, N10154, N1319, N3787);
buf BUF1 (N13502, N13492);
nor NOR4 (N13503, N13500, N5068, N3718, N12938);
and AND2 (N13504, N13503, N8138);
buf BUF1 (N13505, N13478);
or OR2 (N13506, N13486, N5040);
buf BUF1 (N13507, N13496);
buf BUF1 (N13508, N13474);
xor XOR2 (N13509, N13493, N12431);
xor XOR2 (N13510, N13495, N8821);
xor XOR2 (N13511, N13505, N11623);
nor NOR4 (N13512, N13510, N8425, N4308, N6049);
and AND2 (N13513, N13506, N3918);
nor NOR4 (N13514, N13513, N6210, N1767, N359);
nand NAND3 (N13515, N13512, N3826, N2182);
or OR4 (N13516, N13515, N3071, N9480, N9206);
or OR2 (N13517, N13508, N12234);
xor XOR2 (N13518, N13516, N7666);
nand NAND3 (N13519, N13504, N1778, N8698);
or OR2 (N13520, N13511, N12404);
or OR2 (N13521, N13509, N13211);
xor XOR2 (N13522, N13501, N2817);
and AND2 (N13523, N13517, N6350);
or OR2 (N13524, N13519, N5417);
nand NAND4 (N13525, N13523, N2029, N9052, N4659);
or OR2 (N13526, N13518, N5951);
xor XOR2 (N13527, N13524, N6269);
or OR2 (N13528, N13502, N7013);
xor XOR2 (N13529, N13526, N5681);
nor NOR2 (N13530, N13520, N1876);
or OR4 (N13531, N13514, N10838, N2423, N5587);
xor XOR2 (N13532, N13529, N4954);
or OR2 (N13533, N13528, N2867);
not NOT1 (N13534, N13530);
and AND4 (N13535, N13532, N1202, N1354, N4628);
xor XOR2 (N13536, N13522, N11843);
buf BUF1 (N13537, N13525);
xor XOR2 (N13538, N13527, N4199);
buf BUF1 (N13539, N13538);
xor XOR2 (N13540, N13498, N5437);
and AND4 (N13541, N13535, N8576, N11383, N1546);
nand NAND4 (N13542, N13541, N5640, N8961, N11688);
and AND4 (N13543, N13521, N9842, N10350, N9786);
and AND2 (N13544, N13542, N10359);
nand NAND3 (N13545, N13531, N9468, N12946);
xor XOR2 (N13546, N13544, N7885);
or OR2 (N13547, N13546, N2610);
xor XOR2 (N13548, N13534, N3061);
not NOT1 (N13549, N13539);
not NOT1 (N13550, N13533);
nor NOR2 (N13551, N13543, N7465);
buf BUF1 (N13552, N13549);
or OR2 (N13553, N13548, N11207);
xor XOR2 (N13554, N13537, N5492);
not NOT1 (N13555, N13554);
nand NAND3 (N13556, N13507, N769, N6602);
and AND3 (N13557, N13551, N10055, N200);
or OR2 (N13558, N13555, N10743);
buf BUF1 (N13559, N13558);
nor NOR4 (N13560, N13553, N6445, N2325, N10860);
xor XOR2 (N13561, N13559, N4205);
nand NAND2 (N13562, N13545, N1600);
xor XOR2 (N13563, N13562, N7203);
and AND2 (N13564, N13557, N550);
nor NOR3 (N13565, N13547, N11486, N13122);
not NOT1 (N13566, N13540);
xor XOR2 (N13567, N13563, N52);
nor NOR2 (N13568, N13556, N5895);
nor NOR2 (N13569, N13536, N7378);
nor NOR3 (N13570, N13566, N11538, N1085);
and AND2 (N13571, N13565, N2361);
nand NAND4 (N13572, N13571, N8508, N1252, N7503);
buf BUF1 (N13573, N13569);
buf BUF1 (N13574, N13560);
buf BUF1 (N13575, N13561);
xor XOR2 (N13576, N13574, N2269);
or OR2 (N13577, N13575, N10295);
buf BUF1 (N13578, N13572);
buf BUF1 (N13579, N13552);
xor XOR2 (N13580, N13568, N13311);
and AND3 (N13581, N13564, N11507, N12704);
nor NOR3 (N13582, N13570, N12699, N13252);
not NOT1 (N13583, N13576);
nand NAND4 (N13584, N13582, N4960, N10403, N8712);
xor XOR2 (N13585, N13567, N3609);
or OR3 (N13586, N13585, N10825, N8345);
xor XOR2 (N13587, N13577, N10168);
buf BUF1 (N13588, N13579);
and AND2 (N13589, N13584, N2347);
and AND2 (N13590, N13587, N406);
xor XOR2 (N13591, N13590, N6143);
nor NOR3 (N13592, N13583, N7883, N4139);
and AND3 (N13593, N13589, N6141, N1862);
and AND4 (N13594, N13578, N10296, N10217, N8227);
nand NAND2 (N13595, N13592, N1119);
xor XOR2 (N13596, N13581, N4854);
or OR3 (N13597, N13594, N11315, N2590);
not NOT1 (N13598, N13573);
xor XOR2 (N13599, N13580, N12564);
and AND2 (N13600, N13597, N5679);
nand NAND2 (N13601, N13588, N10350);
xor XOR2 (N13602, N13586, N11517);
not NOT1 (N13603, N13601);
nor NOR3 (N13604, N13595, N989, N3380);
and AND3 (N13605, N13599, N10487, N2913);
buf BUF1 (N13606, N13600);
or OR4 (N13607, N13591, N12302, N2727, N12544);
buf BUF1 (N13608, N13598);
not NOT1 (N13609, N13605);
buf BUF1 (N13610, N13608);
not NOT1 (N13611, N13593);
xor XOR2 (N13612, N13610, N8251);
xor XOR2 (N13613, N13602, N12038);
not NOT1 (N13614, N13550);
xor XOR2 (N13615, N13604, N4290);
nor NOR3 (N13616, N13603, N4260, N9013);
not NOT1 (N13617, N13607);
nor NOR2 (N13618, N13616, N1579);
nor NOR2 (N13619, N13606, N12057);
nand NAND2 (N13620, N13609, N3220);
or OR2 (N13621, N13612, N6766);
not NOT1 (N13622, N13611);
and AND4 (N13623, N13615, N352, N13345, N905);
buf BUF1 (N13624, N13621);
nand NAND3 (N13625, N13622, N246, N6187);
and AND3 (N13626, N13596, N4538, N8050);
or OR4 (N13627, N13624, N2505, N780, N1349);
not NOT1 (N13628, N13618);
xor XOR2 (N13629, N13619, N10472);
buf BUF1 (N13630, N13623);
xor XOR2 (N13631, N13614, N10198);
not NOT1 (N13632, N13630);
buf BUF1 (N13633, N13626);
and AND3 (N13634, N13631, N51, N7078);
nand NAND4 (N13635, N13629, N5839, N5916, N4465);
nand NAND2 (N13636, N13617, N6055);
or OR2 (N13637, N13632, N10017);
nor NOR4 (N13638, N13635, N6688, N10420, N13385);
or OR4 (N13639, N13636, N5012, N8892, N9814);
or OR2 (N13640, N13639, N11785);
not NOT1 (N13641, N13620);
and AND3 (N13642, N13634, N9490, N945);
nand NAND2 (N13643, N13638, N5276);
not NOT1 (N13644, N13628);
or OR2 (N13645, N13640, N3463);
not NOT1 (N13646, N13641);
xor XOR2 (N13647, N13613, N8850);
or OR4 (N13648, N13633, N11768, N1059, N13190);
nor NOR3 (N13649, N13644, N12419, N5013);
buf BUF1 (N13650, N13625);
nor NOR3 (N13651, N13646, N2247, N11071);
nor NOR4 (N13652, N13627, N7122, N5920, N11665);
buf BUF1 (N13653, N13650);
nand NAND3 (N13654, N13649, N2374, N4583);
nand NAND2 (N13655, N13654, N1350);
and AND4 (N13656, N13655, N4299, N12153, N5835);
nand NAND3 (N13657, N13656, N9260, N3556);
nand NAND2 (N13658, N13651, N3204);
not NOT1 (N13659, N13657);
nand NAND3 (N13660, N13643, N1892, N4477);
or OR4 (N13661, N13642, N8179, N7863, N9895);
or OR3 (N13662, N13648, N2639, N11053);
not NOT1 (N13663, N13645);
and AND3 (N13664, N13653, N7688, N7724);
or OR3 (N13665, N13637, N11421, N12401);
buf BUF1 (N13666, N13659);
not NOT1 (N13667, N13660);
and AND3 (N13668, N13663, N268, N206);
nor NOR3 (N13669, N13647, N10715, N1230);
not NOT1 (N13670, N13658);
and AND2 (N13671, N13669, N4008);
and AND4 (N13672, N13665, N13299, N3799, N1128);
buf BUF1 (N13673, N13667);
or OR4 (N13674, N13672, N8444, N7548, N11028);
not NOT1 (N13675, N13664);
or OR4 (N13676, N13652, N10860, N11593, N4064);
not NOT1 (N13677, N13673);
buf BUF1 (N13678, N13675);
not NOT1 (N13679, N13666);
not NOT1 (N13680, N13662);
nor NOR3 (N13681, N13677, N9707, N10442);
buf BUF1 (N13682, N13674);
or OR2 (N13683, N13680, N3304);
or OR4 (N13684, N13682, N315, N8516, N8011);
not NOT1 (N13685, N13676);
buf BUF1 (N13686, N13670);
and AND2 (N13687, N13671, N3774);
and AND4 (N13688, N13687, N12590, N7631, N11948);
not NOT1 (N13689, N13684);
not NOT1 (N13690, N13689);
buf BUF1 (N13691, N13685);
and AND4 (N13692, N13686, N3243, N3717, N4155);
not NOT1 (N13693, N13690);
or OR4 (N13694, N13679, N914, N10944, N10033);
or OR2 (N13695, N13681, N2223);
not NOT1 (N13696, N13695);
not NOT1 (N13697, N13691);
buf BUF1 (N13698, N13668);
and AND3 (N13699, N13661, N10668, N10072);
nand NAND3 (N13700, N13696, N7768, N7415);
xor XOR2 (N13701, N13688, N8483);
and AND3 (N13702, N13678, N5557, N6736);
buf BUF1 (N13703, N13701);
or OR4 (N13704, N13683, N13680, N4768, N5618);
nor NOR2 (N13705, N13699, N7909);
and AND3 (N13706, N13703, N4466, N5986);
or OR4 (N13707, N13706, N1055, N11901, N2564);
nand NAND4 (N13708, N13702, N6795, N268, N12081);
buf BUF1 (N13709, N13693);
nand NAND3 (N13710, N13705, N11937, N9560);
buf BUF1 (N13711, N13698);
or OR3 (N13712, N13694, N4016, N6125);
nand NAND4 (N13713, N13707, N12562, N2378, N8667);
or OR3 (N13714, N13709, N9682, N10741);
not NOT1 (N13715, N13697);
nand NAND2 (N13716, N13704, N12180);
or OR4 (N13717, N13710, N1831, N6629, N4221);
nand NAND3 (N13718, N13716, N1191, N11881);
nand NAND2 (N13719, N13718, N4098);
or OR4 (N13720, N13714, N12341, N12096, N11731);
nor NOR3 (N13721, N13719, N9627, N7653);
or OR3 (N13722, N13712, N8521, N8977);
xor XOR2 (N13723, N13711, N7929);
nand NAND2 (N13724, N13715, N4874);
nor NOR3 (N13725, N13700, N5895, N7823);
nand NAND2 (N13726, N13692, N5693);
nor NOR4 (N13727, N13713, N4219, N4553, N8562);
buf BUF1 (N13728, N13724);
buf BUF1 (N13729, N13708);
xor XOR2 (N13730, N13720, N13135);
and AND2 (N13731, N13729, N12333);
nand NAND2 (N13732, N13731, N4475);
nor NOR2 (N13733, N13727, N2538);
or OR4 (N13734, N13728, N13652, N12907, N1300);
nor NOR4 (N13735, N13733, N4370, N10459, N11068);
and AND4 (N13736, N13730, N8056, N10078, N6954);
nand NAND4 (N13737, N13723, N4408, N6358, N4926);
nand NAND3 (N13738, N13721, N214, N9152);
buf BUF1 (N13739, N13732);
buf BUF1 (N13740, N13722);
and AND2 (N13741, N13738, N7415);
not NOT1 (N13742, N13739);
not NOT1 (N13743, N13726);
or OR2 (N13744, N13735, N4827);
or OR4 (N13745, N13725, N8960, N12150, N8531);
nor NOR3 (N13746, N13734, N4843, N6606);
nand NAND2 (N13747, N13741, N7443);
and AND4 (N13748, N13747, N12118, N861, N10178);
xor XOR2 (N13749, N13743, N11312);
not NOT1 (N13750, N13744);
not NOT1 (N13751, N13717);
xor XOR2 (N13752, N13740, N7805);
xor XOR2 (N13753, N13742, N13321);
nand NAND2 (N13754, N13746, N1020);
or OR2 (N13755, N13748, N13580);
buf BUF1 (N13756, N13755);
nand NAND3 (N13757, N13754, N6086, N4581);
nor NOR3 (N13758, N13749, N8360, N13283);
nor NOR4 (N13759, N13752, N9664, N4532, N10678);
or OR2 (N13760, N13753, N9458);
xor XOR2 (N13761, N13757, N13604);
buf BUF1 (N13762, N13756);
nand NAND3 (N13763, N13760, N9485, N3822);
and AND3 (N13764, N13745, N12053, N10226);
nand NAND3 (N13765, N13759, N6787, N1428);
buf BUF1 (N13766, N13750);
xor XOR2 (N13767, N13736, N793);
or OR2 (N13768, N13761, N6942);
and AND3 (N13769, N13758, N1631, N11254);
nand NAND3 (N13770, N13766, N10870, N11418);
nand NAND4 (N13771, N13762, N2608, N965, N9381);
nand NAND4 (N13772, N13770, N12086, N8274, N2621);
xor XOR2 (N13773, N13767, N7909);
buf BUF1 (N13774, N13764);
nor NOR3 (N13775, N13768, N3802, N9152);
and AND4 (N13776, N13772, N13043, N5290, N11096);
buf BUF1 (N13777, N13771);
or OR2 (N13778, N13777, N10381);
nand NAND3 (N13779, N13751, N12056, N408);
nor NOR2 (N13780, N13779, N2425);
buf BUF1 (N13781, N13776);
and AND3 (N13782, N13780, N2345, N2995);
not NOT1 (N13783, N13763);
or OR2 (N13784, N13782, N2657);
or OR4 (N13785, N13774, N8253, N10799, N11364);
not NOT1 (N13786, N13773);
not NOT1 (N13787, N13778);
and AND2 (N13788, N13786, N9019);
nand NAND2 (N13789, N13785, N6111);
nand NAND3 (N13790, N13784, N10686, N6111);
and AND3 (N13791, N13788, N9906, N4887);
nor NOR3 (N13792, N13789, N5759, N2811);
xor XOR2 (N13793, N13737, N4452);
and AND2 (N13794, N13791, N5324);
xor XOR2 (N13795, N13787, N3355);
buf BUF1 (N13796, N13795);
buf BUF1 (N13797, N13765);
buf BUF1 (N13798, N13781);
or OR4 (N13799, N13792, N11498, N1270, N7816);
not NOT1 (N13800, N13796);
or OR3 (N13801, N13800, N2384, N5068);
or OR2 (N13802, N13775, N1315);
buf BUF1 (N13803, N13799);
nor NOR3 (N13804, N13794, N8380, N5239);
or OR2 (N13805, N13793, N1690);
nor NOR2 (N13806, N13804, N8206);
nor NOR2 (N13807, N13783, N8855);
and AND3 (N13808, N13797, N1711, N9889);
and AND3 (N13809, N13802, N349, N11286);
and AND3 (N13810, N13806, N8266, N8316);
nor NOR3 (N13811, N13803, N3663, N4445);
buf BUF1 (N13812, N13801);
not NOT1 (N13813, N13798);
or OR3 (N13814, N13790, N7053, N9065);
or OR4 (N13815, N13813, N8343, N13797, N6194);
xor XOR2 (N13816, N13810, N2476);
nor NOR4 (N13817, N13807, N9764, N222, N3774);
xor XOR2 (N13818, N13815, N3845);
or OR2 (N13819, N13814, N1720);
and AND4 (N13820, N13809, N6512, N13733, N56);
nor NOR2 (N13821, N13817, N9707);
or OR2 (N13822, N13816, N4477);
and AND2 (N13823, N13820, N1446);
nor NOR2 (N13824, N13819, N6847);
or OR3 (N13825, N13808, N9457, N6546);
xor XOR2 (N13826, N13812, N13464);
not NOT1 (N13827, N13823);
nor NOR2 (N13828, N13824, N3531);
xor XOR2 (N13829, N13818, N2351);
and AND4 (N13830, N13826, N7079, N12450, N6218);
and AND4 (N13831, N13829, N8055, N2658, N3446);
xor XOR2 (N13832, N13828, N3864);
or OR3 (N13833, N13827, N12545, N1688);
not NOT1 (N13834, N13822);
or OR3 (N13835, N13830, N4618, N8074);
or OR3 (N13836, N13832, N3588, N10529);
xor XOR2 (N13837, N13825, N2698);
and AND2 (N13838, N13821, N5007);
nor NOR2 (N13839, N13835, N2029);
and AND2 (N13840, N13833, N8913);
not NOT1 (N13841, N13811);
or OR3 (N13842, N13840, N4773, N7801);
nor NOR4 (N13843, N13837, N3171, N4147, N5157);
xor XOR2 (N13844, N13831, N2378);
nor NOR3 (N13845, N13839, N6371, N6741);
xor XOR2 (N13846, N13805, N9538);
xor XOR2 (N13847, N13838, N2913);
nand NAND4 (N13848, N13843, N3617, N3173, N13218);
buf BUF1 (N13849, N13847);
not NOT1 (N13850, N13844);
xor XOR2 (N13851, N13848, N5345);
and AND2 (N13852, N13849, N2804);
nand NAND2 (N13853, N13836, N3139);
and AND4 (N13854, N13841, N8120, N13394, N5087);
and AND4 (N13855, N13769, N1487, N13779, N10120);
buf BUF1 (N13856, N13846);
nand NAND3 (N13857, N13853, N12775, N558);
nor NOR4 (N13858, N13852, N5891, N13414, N5494);
nand NAND3 (N13859, N13842, N585, N10722);
not NOT1 (N13860, N13845);
or OR4 (N13861, N13857, N5468, N11461, N5133);
not NOT1 (N13862, N13861);
buf BUF1 (N13863, N13834);
xor XOR2 (N13864, N13860, N1188);
buf BUF1 (N13865, N13850);
nor NOR4 (N13866, N13859, N7403, N9273, N3538);
nand NAND3 (N13867, N13851, N275, N8173);
nor NOR2 (N13868, N13867, N13321);
and AND4 (N13869, N13858, N9596, N10748, N6320);
nand NAND4 (N13870, N13869, N6518, N8044, N3405);
not NOT1 (N13871, N13866);
not NOT1 (N13872, N13863);
buf BUF1 (N13873, N13862);
or OR2 (N13874, N13868, N13355);
buf BUF1 (N13875, N13865);
nand NAND2 (N13876, N13870, N5089);
buf BUF1 (N13877, N13874);
nand NAND2 (N13878, N13873, N2802);
nor NOR4 (N13879, N13872, N10280, N7050, N8813);
buf BUF1 (N13880, N13877);
and AND3 (N13881, N13856, N6154, N5322);
not NOT1 (N13882, N13879);
nor NOR2 (N13883, N13875, N1071);
not NOT1 (N13884, N13871);
xor XOR2 (N13885, N13855, N1544);
xor XOR2 (N13886, N13864, N12710);
buf BUF1 (N13887, N13878);
and AND3 (N13888, N13881, N11260, N7696);
and AND4 (N13889, N13886, N13598, N10471, N3237);
nand NAND3 (N13890, N13880, N10554, N6055);
not NOT1 (N13891, N13882);
xor XOR2 (N13892, N13854, N4841);
xor XOR2 (N13893, N13885, N1103);
nor NOR2 (N13894, N13883, N2197);
buf BUF1 (N13895, N13891);
and AND2 (N13896, N13889, N2782);
nand NAND2 (N13897, N13892, N11962);
or OR3 (N13898, N13876, N10688, N10759);
or OR3 (N13899, N13890, N4877, N2159);
nor NOR2 (N13900, N13894, N10940);
or OR4 (N13901, N13884, N1782, N12966, N9322);
not NOT1 (N13902, N13899);
and AND4 (N13903, N13902, N353, N10820, N12335);
xor XOR2 (N13904, N13895, N11259);
xor XOR2 (N13905, N13888, N6476);
xor XOR2 (N13906, N13896, N11779);
not NOT1 (N13907, N13887);
nand NAND4 (N13908, N13901, N10224, N1885, N9004);
nand NAND3 (N13909, N13904, N9688, N191);
not NOT1 (N13910, N13907);
or OR2 (N13911, N13909, N3300);
nor NOR4 (N13912, N13910, N10036, N7626, N2541);
buf BUF1 (N13913, N13908);
or OR3 (N13914, N13897, N13719, N12926);
and AND2 (N13915, N13911, N173);
xor XOR2 (N13916, N13905, N5392);
not NOT1 (N13917, N13898);
or OR4 (N13918, N13893, N10575, N6020, N4697);
nand NAND3 (N13919, N13913, N74, N5856);
xor XOR2 (N13920, N13918, N12108);
not NOT1 (N13921, N13903);
and AND4 (N13922, N13916, N12142, N7026, N6068);
xor XOR2 (N13923, N13914, N4747);
and AND3 (N13924, N13922, N9938, N10109);
nor NOR3 (N13925, N13906, N6269, N5822);
not NOT1 (N13926, N13912);
and AND4 (N13927, N13923, N5152, N13571, N1746);
nor NOR2 (N13928, N13915, N1101);
not NOT1 (N13929, N13927);
xor XOR2 (N13930, N13917, N11060);
xor XOR2 (N13931, N13926, N6782);
or OR3 (N13932, N13930, N8570, N13182);
and AND3 (N13933, N13932, N13797, N592);
and AND2 (N13934, N13920, N3569);
buf BUF1 (N13935, N13929);
buf BUF1 (N13936, N13900);
not NOT1 (N13937, N13924);
or OR3 (N13938, N13921, N2413, N5661);
and AND2 (N13939, N13931, N1408);
and AND2 (N13940, N13935, N7565);
not NOT1 (N13941, N13934);
xor XOR2 (N13942, N13940, N4154);
not NOT1 (N13943, N13938);
buf BUF1 (N13944, N13941);
or OR2 (N13945, N13939, N12476);
xor XOR2 (N13946, N13928, N3880);
buf BUF1 (N13947, N13919);
or OR3 (N13948, N13933, N2103, N9490);
or OR2 (N13949, N13936, N9675);
nor NOR2 (N13950, N13947, N6307);
and AND3 (N13951, N13950, N2308, N9214);
or OR2 (N13952, N13945, N7849);
and AND4 (N13953, N13943, N7677, N2682, N4433);
buf BUF1 (N13954, N13937);
buf BUF1 (N13955, N13946);
and AND3 (N13956, N13942, N13216, N1657);
nor NOR2 (N13957, N13952, N2135);
nand NAND2 (N13958, N13951, N6962);
nor NOR2 (N13959, N13957, N10710);
buf BUF1 (N13960, N13948);
and AND2 (N13961, N13958, N8852);
and AND3 (N13962, N13953, N4840, N11555);
nand NAND2 (N13963, N13956, N9864);
nand NAND2 (N13964, N13963, N2187);
nand NAND3 (N13965, N13955, N6315, N5918);
and AND2 (N13966, N13959, N8075);
and AND4 (N13967, N13962, N430, N13414, N4628);
nor NOR3 (N13968, N13965, N2724, N8245);
nand NAND4 (N13969, N13960, N10966, N8867, N13065);
nand NAND3 (N13970, N13969, N12466, N13822);
or OR2 (N13971, N13944, N9084);
or OR3 (N13972, N13966, N152, N4992);
nand NAND4 (N13973, N13972, N4496, N1121, N11820);
not NOT1 (N13974, N13961);
and AND4 (N13975, N13971, N7557, N6770, N626);
xor XOR2 (N13976, N13954, N2776);
nand NAND2 (N13977, N13967, N3149);
not NOT1 (N13978, N13949);
nand NAND2 (N13979, N13968, N7959);
and AND4 (N13980, N13978, N10587, N10410, N8966);
buf BUF1 (N13981, N13979);
nor NOR4 (N13982, N13974, N13408, N10911, N7779);
nor NOR4 (N13983, N13973, N2389, N11795, N10749);
not NOT1 (N13984, N13980);
xor XOR2 (N13985, N13970, N7293);
nand NAND2 (N13986, N13981, N1538);
or OR3 (N13987, N13975, N12889, N1837);
not NOT1 (N13988, N13986);
and AND4 (N13989, N13983, N9981, N178, N10689);
buf BUF1 (N13990, N13989);
xor XOR2 (N13991, N13988, N4913);
and AND3 (N13992, N13985, N8695, N4141);
buf BUF1 (N13993, N13925);
or OR2 (N13994, N13990, N3967);
nand NAND3 (N13995, N13994, N7024, N12028);
not NOT1 (N13996, N13993);
or OR4 (N13997, N13964, N9368, N10331, N2482);
xor XOR2 (N13998, N13991, N4860);
or OR4 (N13999, N13982, N5927, N33, N10189);
buf BUF1 (N14000, N13995);
xor XOR2 (N14001, N13996, N1709);
xor XOR2 (N14002, N13998, N1228);
not NOT1 (N14003, N13987);
nor NOR3 (N14004, N13984, N7417, N10056);
nand NAND2 (N14005, N13977, N12303);
xor XOR2 (N14006, N14001, N3255);
nand NAND3 (N14007, N14002, N13929, N3634);
not NOT1 (N14008, N14000);
and AND3 (N14009, N13992, N2618, N3107);
or OR3 (N14010, N14004, N2142, N8474);
or OR4 (N14011, N14006, N7538, N8557, N1082);
and AND2 (N14012, N13997, N12566);
or OR2 (N14013, N14008, N4635);
and AND2 (N14014, N14009, N7672);
xor XOR2 (N14015, N13976, N7038);
and AND4 (N14016, N14010, N3053, N8838, N6661);
not NOT1 (N14017, N14015);
xor XOR2 (N14018, N14012, N9978);
nand NAND2 (N14019, N14018, N6206);
nor NOR3 (N14020, N14017, N7465, N2092);
buf BUF1 (N14021, N14003);
nand NAND4 (N14022, N14011, N4797, N10800, N5927);
buf BUF1 (N14023, N14014);
nand NAND4 (N14024, N13999, N1517, N336, N6941);
or OR2 (N14025, N14020, N11520);
and AND3 (N14026, N14013, N11787, N9104);
xor XOR2 (N14027, N14024, N6017);
nor NOR2 (N14028, N14016, N4128);
nor NOR4 (N14029, N14021, N12667, N8055, N11598);
xor XOR2 (N14030, N14022, N8111);
xor XOR2 (N14031, N14005, N11159);
not NOT1 (N14032, N14027);
nor NOR4 (N14033, N14007, N8223, N460, N9778);
nor NOR2 (N14034, N14031, N8722);
nor NOR2 (N14035, N14026, N1207);
buf BUF1 (N14036, N14019);
and AND4 (N14037, N14034, N2879, N3265, N3846);
or OR4 (N14038, N14036, N679, N7743, N2665);
not NOT1 (N14039, N14038);
or OR4 (N14040, N14030, N1341, N7681, N5340);
and AND3 (N14041, N14037, N7677, N498);
or OR2 (N14042, N14028, N13711);
and AND4 (N14043, N14039, N2420, N6742, N10797);
nand NAND3 (N14044, N14041, N12756, N1687);
xor XOR2 (N14045, N14044, N12353);
or OR3 (N14046, N14023, N11765, N6323);
buf BUF1 (N14047, N14042);
buf BUF1 (N14048, N14046);
nand NAND2 (N14049, N14033, N4429);
buf BUF1 (N14050, N14035);
buf BUF1 (N14051, N14049);
or OR3 (N14052, N14032, N9263, N4050);
and AND4 (N14053, N14040, N9929, N6506, N10975);
or OR2 (N14054, N14045, N4826);
buf BUF1 (N14055, N14029);
and AND4 (N14056, N14043, N12917, N3234, N4819);
xor XOR2 (N14057, N14050, N1450);
not NOT1 (N14058, N14053);
or OR3 (N14059, N14048, N8719, N11956);
and AND4 (N14060, N14025, N5705, N11713, N9419);
and AND4 (N14061, N14059, N13329, N5420, N6394);
nor NOR2 (N14062, N14060, N10949);
nand NAND4 (N14063, N14052, N9743, N2199, N12861);
xor XOR2 (N14064, N14063, N8904);
or OR3 (N14065, N14047, N569, N13894);
not NOT1 (N14066, N14062);
or OR4 (N14067, N14051, N12477, N719, N7269);
and AND2 (N14068, N14065, N8646);
nand NAND4 (N14069, N14054, N7472, N4295, N13959);
and AND2 (N14070, N14056, N3548);
nor NOR4 (N14071, N14061, N6960, N10765, N3899);
xor XOR2 (N14072, N14066, N1798);
and AND4 (N14073, N14068, N5444, N1565, N13418);
nor NOR4 (N14074, N14058, N10358, N4657, N5878);
xor XOR2 (N14075, N14069, N8476);
nor NOR4 (N14076, N14057, N11008, N4487, N2542);
or OR2 (N14077, N14070, N3477);
nor NOR2 (N14078, N14076, N7220);
not NOT1 (N14079, N14077);
buf BUF1 (N14080, N14079);
not NOT1 (N14081, N14071);
not NOT1 (N14082, N14078);
nand NAND2 (N14083, N14072, N6882);
not NOT1 (N14084, N14074);
or OR2 (N14085, N14064, N11966);
xor XOR2 (N14086, N14084, N6259);
nand NAND3 (N14087, N14075, N8388, N5707);
not NOT1 (N14088, N14067);
nor NOR4 (N14089, N14086, N11959, N9648, N3916);
nand NAND4 (N14090, N14082, N2127, N12723, N10373);
nand NAND4 (N14091, N14090, N1128, N3931, N6154);
xor XOR2 (N14092, N14080, N4482);
not NOT1 (N14093, N14083);
xor XOR2 (N14094, N14092, N380);
not NOT1 (N14095, N14093);
nor NOR2 (N14096, N14055, N10249);
not NOT1 (N14097, N14081);
nor NOR2 (N14098, N14091, N6216);
or OR3 (N14099, N14088, N3743, N7754);
nand NAND4 (N14100, N14098, N12633, N1377, N4403);
xor XOR2 (N14101, N14096, N11649);
and AND3 (N14102, N14073, N3025, N6589);
not NOT1 (N14103, N14085);
nor NOR3 (N14104, N14094, N200, N10789);
not NOT1 (N14105, N14095);
buf BUF1 (N14106, N14102);
buf BUF1 (N14107, N14097);
buf BUF1 (N14108, N14087);
not NOT1 (N14109, N14105);
xor XOR2 (N14110, N14106, N9011);
buf BUF1 (N14111, N14103);
xor XOR2 (N14112, N14108, N1393);
not NOT1 (N14113, N14100);
not NOT1 (N14114, N14109);
buf BUF1 (N14115, N14111);
and AND4 (N14116, N14112, N3387, N2398, N12855);
and AND3 (N14117, N14110, N10380, N13002);
or OR4 (N14118, N14117, N12263, N4697, N5169);
or OR2 (N14119, N14114, N6647);
xor XOR2 (N14120, N14101, N6417);
buf BUF1 (N14121, N14119);
nand NAND3 (N14122, N14107, N9066, N12954);
not NOT1 (N14123, N14089);
and AND2 (N14124, N14099, N2442);
xor XOR2 (N14125, N14120, N8498);
not NOT1 (N14126, N14113);
not NOT1 (N14127, N14104);
or OR3 (N14128, N14122, N525, N1963);
nand NAND4 (N14129, N14116, N12722, N10710, N8151);
xor XOR2 (N14130, N14115, N13835);
not NOT1 (N14131, N14123);
xor XOR2 (N14132, N14127, N8647);
buf BUF1 (N14133, N14132);
and AND2 (N14134, N14130, N13764);
and AND3 (N14135, N14131, N13734, N7619);
nor NOR2 (N14136, N14129, N69);
buf BUF1 (N14137, N14128);
or OR3 (N14138, N14121, N13589, N4773);
buf BUF1 (N14139, N14118);
nor NOR3 (N14140, N14125, N3884, N1295);
and AND4 (N14141, N14135, N2374, N2613, N7911);
nor NOR4 (N14142, N14124, N13522, N12007, N5849);
nor NOR4 (N14143, N14134, N8107, N13982, N12847);
nor NOR3 (N14144, N14141, N10735, N5370);
not NOT1 (N14145, N14126);
and AND3 (N14146, N14138, N13259, N8304);
not NOT1 (N14147, N14136);
buf BUF1 (N14148, N14133);
and AND3 (N14149, N14145, N757, N2808);
not NOT1 (N14150, N14148);
nor NOR4 (N14151, N14147, N7151, N13681, N2469);
and AND3 (N14152, N14139, N5695, N6127);
xor XOR2 (N14153, N14150, N977);
or OR4 (N14154, N14140, N5589, N9704, N4910);
and AND4 (N14155, N14153, N13478, N13389, N10546);
and AND2 (N14156, N14144, N6365);
not NOT1 (N14157, N14155);
xor XOR2 (N14158, N14156, N12071);
nor NOR4 (N14159, N14158, N3161, N4997, N11875);
xor XOR2 (N14160, N14137, N4904);
nor NOR3 (N14161, N14146, N6895, N10217);
buf BUF1 (N14162, N14142);
and AND3 (N14163, N14149, N11467, N2999);
xor XOR2 (N14164, N14152, N3787);
xor XOR2 (N14165, N14151, N4538);
not NOT1 (N14166, N14159);
xor XOR2 (N14167, N14161, N7461);
and AND4 (N14168, N14160, N11262, N8192, N3562);
not NOT1 (N14169, N14165);
nor NOR2 (N14170, N14166, N8264);
or OR3 (N14171, N14157, N11845, N12436);
buf BUF1 (N14172, N14171);
xor XOR2 (N14173, N14143, N1369);
or OR4 (N14174, N14170, N5072, N5670, N4043);
not NOT1 (N14175, N14173);
xor XOR2 (N14176, N14172, N11441);
nand NAND4 (N14177, N14163, N4312, N2964, N5369);
nand NAND4 (N14178, N14176, N6232, N3450, N7778);
or OR4 (N14179, N14168, N6192, N11944, N4245);
not NOT1 (N14180, N14169);
or OR4 (N14181, N14167, N1256, N382, N2214);
and AND2 (N14182, N14179, N8330);
and AND3 (N14183, N14174, N5715, N3814);
or OR3 (N14184, N14178, N9948, N1519);
nor NOR2 (N14185, N14175, N11035);
nor NOR2 (N14186, N14185, N7811);
or OR2 (N14187, N14184, N11495);
nand NAND2 (N14188, N14182, N953);
and AND4 (N14189, N14183, N8192, N9941, N604);
nor NOR2 (N14190, N14177, N12150);
not NOT1 (N14191, N14190);
nand NAND4 (N14192, N14180, N5809, N3965, N11123);
nor NOR3 (N14193, N14186, N1447, N9167);
nand NAND3 (N14194, N14162, N2032, N836);
or OR4 (N14195, N14181, N4404, N9706, N5427);
not NOT1 (N14196, N14193);
xor XOR2 (N14197, N14191, N12994);
xor XOR2 (N14198, N14194, N4747);
nand NAND4 (N14199, N14154, N1144, N4742, N2481);
and AND2 (N14200, N14198, N2587);
and AND4 (N14201, N14196, N6791, N9075, N3648);
nor NOR3 (N14202, N14192, N7194, N3494);
not NOT1 (N14203, N14195);
nand NAND3 (N14204, N14189, N14073, N12695);
not NOT1 (N14205, N14200);
xor XOR2 (N14206, N14188, N3046);
or OR4 (N14207, N14202, N768, N1081, N1661);
buf BUF1 (N14208, N14197);
buf BUF1 (N14209, N14207);
nor NOR2 (N14210, N14203, N3377);
or OR4 (N14211, N14201, N11477, N2587, N4948);
and AND2 (N14212, N14211, N5572);
and AND4 (N14213, N14212, N50, N9749, N13242);
nor NOR4 (N14214, N14209, N4821, N3519, N10858);
xor XOR2 (N14215, N14210, N9890);
and AND3 (N14216, N14213, N13970, N5776);
xor XOR2 (N14217, N14208, N4216);
xor XOR2 (N14218, N14217, N917);
and AND3 (N14219, N14164, N4480, N2825);
xor XOR2 (N14220, N14216, N14007);
or OR2 (N14221, N14219, N14016);
and AND4 (N14222, N14218, N2482, N13148, N12595);
nor NOR2 (N14223, N14221, N8020);
not NOT1 (N14224, N14214);
nand NAND4 (N14225, N14206, N11813, N643, N3134);
nor NOR3 (N14226, N14225, N1216, N4921);
or OR2 (N14227, N14224, N11606);
or OR3 (N14228, N14204, N2665, N6488);
or OR4 (N14229, N14222, N10568, N7723, N9790);
nand NAND3 (N14230, N14228, N11884, N7867);
or OR4 (N14231, N14187, N4666, N10107, N7476);
nor NOR4 (N14232, N14230, N6883, N10380, N13435);
not NOT1 (N14233, N14205);
nor NOR3 (N14234, N14199, N280, N6665);
not NOT1 (N14235, N14234);
nor NOR3 (N14236, N14220, N867, N2912);
nor NOR3 (N14237, N14236, N7373, N1253);
not NOT1 (N14238, N14231);
nor NOR2 (N14239, N14226, N2890);
xor XOR2 (N14240, N14232, N4691);
nand NAND3 (N14241, N14215, N3612, N5354);
xor XOR2 (N14242, N14235, N7255);
not NOT1 (N14243, N14239);
or OR2 (N14244, N14233, N11611);
not NOT1 (N14245, N14242);
not NOT1 (N14246, N14227);
nand NAND2 (N14247, N14243, N11523);
and AND4 (N14248, N14238, N8119, N8255, N4940);
and AND4 (N14249, N14246, N10834, N9937, N1979);
and AND4 (N14250, N14240, N3569, N4432, N8335);
buf BUF1 (N14251, N14229);
nand NAND4 (N14252, N14247, N3167, N9004, N13207);
buf BUF1 (N14253, N14248);
xor XOR2 (N14254, N14252, N3777);
and AND4 (N14255, N14251, N10227, N12168, N1094);
buf BUF1 (N14256, N14253);
or OR4 (N14257, N14223, N12816, N9497, N11290);
or OR3 (N14258, N14250, N228, N8835);
nand NAND4 (N14259, N14237, N5171, N2030, N13280);
buf BUF1 (N14260, N14259);
or OR3 (N14261, N14257, N11638, N11672);
or OR2 (N14262, N14241, N4395);
or OR2 (N14263, N14244, N6749);
not NOT1 (N14264, N14258);
not NOT1 (N14265, N14254);
and AND2 (N14266, N14261, N14149);
nor NOR2 (N14267, N14260, N9880);
buf BUF1 (N14268, N14249);
buf BUF1 (N14269, N14268);
xor XOR2 (N14270, N14265, N1375);
or OR4 (N14271, N14270, N13362, N10036, N11058);
buf BUF1 (N14272, N14263);
or OR2 (N14273, N14266, N12822);
not NOT1 (N14274, N14262);
not NOT1 (N14275, N14273);
not NOT1 (N14276, N14272);
and AND3 (N14277, N14264, N1808, N13869);
or OR3 (N14278, N14269, N6519, N3710);
or OR3 (N14279, N14276, N664, N7999);
and AND3 (N14280, N14274, N4859, N7366);
or OR2 (N14281, N14255, N7376);
nor NOR4 (N14282, N14281, N1310, N9193, N7219);
buf BUF1 (N14283, N14271);
and AND2 (N14284, N14280, N10596);
nor NOR2 (N14285, N14279, N10741);
not NOT1 (N14286, N14275);
or OR4 (N14287, N14277, N620, N11580, N7730);
xor XOR2 (N14288, N14256, N3932);
buf BUF1 (N14289, N14278);
buf BUF1 (N14290, N14288);
buf BUF1 (N14291, N14284);
or OR2 (N14292, N14245, N12468);
xor XOR2 (N14293, N14285, N6443);
nand NAND3 (N14294, N14287, N939, N601);
nand NAND2 (N14295, N14267, N5469);
xor XOR2 (N14296, N14283, N13066);
buf BUF1 (N14297, N14296);
nor NOR2 (N14298, N14295, N5297);
xor XOR2 (N14299, N14292, N1717);
or OR2 (N14300, N14282, N9205);
nand NAND3 (N14301, N14293, N2672, N3595);
not NOT1 (N14302, N14298);
xor XOR2 (N14303, N14294, N1851);
and AND3 (N14304, N14301, N6680, N4503);
not NOT1 (N14305, N14286);
xor XOR2 (N14306, N14302, N12220);
or OR2 (N14307, N14299, N1849);
and AND3 (N14308, N14291, N2514, N4205);
or OR2 (N14309, N14307, N12984);
and AND3 (N14310, N14309, N5619, N6265);
buf BUF1 (N14311, N14297);
nand NAND4 (N14312, N14305, N6958, N10434, N5857);
not NOT1 (N14313, N14306);
buf BUF1 (N14314, N14312);
or OR4 (N14315, N14313, N5827, N12430, N2144);
nor NOR3 (N14316, N14303, N3663, N3929);
not NOT1 (N14317, N14308);
xor XOR2 (N14318, N14315, N3495);
or OR4 (N14319, N14318, N273, N483, N10306);
nand NAND2 (N14320, N14311, N4007);
nor NOR3 (N14321, N14300, N6986, N7557);
nand NAND4 (N14322, N14319, N7731, N9787, N9102);
buf BUF1 (N14323, N14316);
not NOT1 (N14324, N14314);
buf BUF1 (N14325, N14289);
nor NOR2 (N14326, N14322, N9294);
not NOT1 (N14327, N14290);
and AND4 (N14328, N14327, N12449, N5380, N1220);
and AND4 (N14329, N14310, N4765, N2473, N7483);
and AND2 (N14330, N14324, N12728);
buf BUF1 (N14331, N14304);
xor XOR2 (N14332, N14325, N6558);
buf BUF1 (N14333, N14328);
or OR2 (N14334, N14326, N7974);
nand NAND3 (N14335, N14320, N1982, N11417);
not NOT1 (N14336, N14329);
buf BUF1 (N14337, N14317);
buf BUF1 (N14338, N14335);
or OR3 (N14339, N14338, N1582, N11745);
not NOT1 (N14340, N14321);
buf BUF1 (N14341, N14331);
xor XOR2 (N14342, N14334, N13082);
nor NOR2 (N14343, N14340, N1022);
and AND4 (N14344, N14341, N4598, N5386, N11187);
or OR4 (N14345, N14343, N12399, N10047, N8809);
or OR2 (N14346, N14332, N14034);
not NOT1 (N14347, N14330);
not NOT1 (N14348, N14345);
buf BUF1 (N14349, N14333);
or OR2 (N14350, N14344, N10835);
and AND2 (N14351, N14339, N9451);
not NOT1 (N14352, N14348);
or OR4 (N14353, N14349, N4967, N6332, N12694);
nor NOR3 (N14354, N14353, N13519, N4854);
or OR2 (N14355, N14323, N13259);
and AND4 (N14356, N14350, N12952, N7545, N2778);
nor NOR4 (N14357, N14356, N14143, N5306, N5991);
or OR2 (N14358, N14352, N8559);
nand NAND2 (N14359, N14355, N5158);
and AND2 (N14360, N14347, N9735);
not NOT1 (N14361, N14358);
not NOT1 (N14362, N14346);
nor NOR2 (N14363, N14351, N12558);
or OR2 (N14364, N14336, N3886);
nand NAND3 (N14365, N14342, N6762, N9071);
and AND4 (N14366, N14361, N13623, N12308, N5808);
buf BUF1 (N14367, N14357);
or OR2 (N14368, N14359, N7982);
nor NOR4 (N14369, N14367, N2379, N7229, N5635);
not NOT1 (N14370, N14369);
not NOT1 (N14371, N14368);
nor NOR3 (N14372, N14362, N4616, N7328);
nand NAND4 (N14373, N14337, N10282, N9640, N1186);
nor NOR4 (N14374, N14360, N4899, N12004, N6076);
xor XOR2 (N14375, N14373, N8789);
xor XOR2 (N14376, N14365, N12197);
and AND3 (N14377, N14370, N5485, N4962);
buf BUF1 (N14378, N14366);
not NOT1 (N14379, N14376);
nand NAND3 (N14380, N14354, N9300, N3462);
buf BUF1 (N14381, N14377);
xor XOR2 (N14382, N14364, N14269);
or OR4 (N14383, N14372, N2132, N8512, N14055);
and AND4 (N14384, N14381, N7447, N5497, N13882);
buf BUF1 (N14385, N14374);
nor NOR4 (N14386, N14382, N5173, N10455, N1113);
xor XOR2 (N14387, N14380, N6557);
xor XOR2 (N14388, N14387, N2201);
and AND2 (N14389, N14363, N7362);
nand NAND3 (N14390, N14389, N7483, N190);
nor NOR2 (N14391, N14375, N14157);
not NOT1 (N14392, N14386);
or OR2 (N14393, N14388, N13377);
buf BUF1 (N14394, N14391);
nor NOR2 (N14395, N14394, N1517);
not NOT1 (N14396, N14385);
or OR3 (N14397, N14371, N8017, N5118);
nand NAND3 (N14398, N14384, N10857, N11379);
xor XOR2 (N14399, N14397, N6879);
nand NAND2 (N14400, N14396, N13086);
and AND3 (N14401, N14399, N12883, N10539);
buf BUF1 (N14402, N14378);
nor NOR3 (N14403, N14392, N5597, N4390);
not NOT1 (N14404, N14393);
and AND3 (N14405, N14383, N10300, N1214);
not NOT1 (N14406, N14390);
and AND2 (N14407, N14379, N11019);
xor XOR2 (N14408, N14398, N662);
xor XOR2 (N14409, N14405, N9079);
nor NOR4 (N14410, N14402, N8312, N12708, N6612);
nor NOR3 (N14411, N14395, N13327, N3623);
xor XOR2 (N14412, N14408, N159);
and AND3 (N14413, N14411, N1398, N7301);
and AND2 (N14414, N14401, N5832);
or OR4 (N14415, N14404, N361, N4304, N8593);
xor XOR2 (N14416, N14410, N6722);
not NOT1 (N14417, N14416);
not NOT1 (N14418, N14413);
nor NOR4 (N14419, N14403, N3944, N6006, N11448);
or OR4 (N14420, N14419, N2802, N12538, N11410);
nand NAND2 (N14421, N14406, N8327);
and AND4 (N14422, N14412, N467, N12529, N1021);
buf BUF1 (N14423, N14418);
nor NOR3 (N14424, N14407, N6914, N12785);
nor NOR4 (N14425, N14423, N2370, N10924, N12979);
xor XOR2 (N14426, N14424, N10308);
and AND3 (N14427, N14409, N9174, N6410);
xor XOR2 (N14428, N14417, N8389);
not NOT1 (N14429, N14414);
xor XOR2 (N14430, N14427, N6995);
nor NOR3 (N14431, N14429, N13182, N6036);
not NOT1 (N14432, N14415);
not NOT1 (N14433, N14425);
or OR3 (N14434, N14422, N7759, N5744);
xor XOR2 (N14435, N14432, N9930);
nor NOR4 (N14436, N14428, N4376, N10313, N7801);
and AND4 (N14437, N14421, N4092, N6440, N5335);
or OR2 (N14438, N14433, N9934);
buf BUF1 (N14439, N14438);
nand NAND2 (N14440, N14434, N7772);
buf BUF1 (N14441, N14431);
not NOT1 (N14442, N14400);
and AND3 (N14443, N14437, N12960, N8878);
not NOT1 (N14444, N14443);
nand NAND2 (N14445, N14436, N9279);
nand NAND2 (N14446, N14426, N14031);
not NOT1 (N14447, N14430);
or OR2 (N14448, N14445, N5168);
or OR3 (N14449, N14448, N9047, N7416);
xor XOR2 (N14450, N14442, N4995);
nor NOR2 (N14451, N14446, N6442);
nand NAND2 (N14452, N14444, N13674);
and AND2 (N14453, N14451, N3291);
nand NAND3 (N14454, N14453, N3395, N12655);
buf BUF1 (N14455, N14452);
not NOT1 (N14456, N14439);
xor XOR2 (N14457, N14441, N3294);
and AND2 (N14458, N14449, N9223);
buf BUF1 (N14459, N14420);
buf BUF1 (N14460, N14455);
or OR2 (N14461, N14457, N9738);
buf BUF1 (N14462, N14461);
nor NOR4 (N14463, N14440, N9279, N2832, N11370);
not NOT1 (N14464, N14450);
not NOT1 (N14465, N14462);
xor XOR2 (N14466, N14435, N12238);
nand NAND2 (N14467, N14463, N6609);
or OR2 (N14468, N14467, N8756);
or OR2 (N14469, N14458, N5264);
nand NAND4 (N14470, N14459, N12002, N12499, N7840);
or OR4 (N14471, N14468, N8905, N8342, N10917);
and AND2 (N14472, N14470, N10224);
or OR3 (N14473, N14460, N2998, N3337);
nor NOR2 (N14474, N14454, N11092);
not NOT1 (N14475, N14472);
xor XOR2 (N14476, N14447, N9381);
nand NAND3 (N14477, N14464, N9181, N2931);
nand NAND4 (N14478, N14465, N5957, N4133, N3044);
and AND3 (N14479, N14473, N6432, N5643);
nor NOR3 (N14480, N14479, N9742, N2196);
or OR3 (N14481, N14474, N8506, N11756);
xor XOR2 (N14482, N14469, N2269);
not NOT1 (N14483, N14456);
not NOT1 (N14484, N14477);
xor XOR2 (N14485, N14482, N4043);
nand NAND3 (N14486, N14483, N5924, N4153);
and AND3 (N14487, N14480, N455, N9723);
not NOT1 (N14488, N14471);
buf BUF1 (N14489, N14475);
nand NAND4 (N14490, N14488, N1898, N2562, N8009);
xor XOR2 (N14491, N14489, N3905);
nand NAND3 (N14492, N14476, N892, N5527);
not NOT1 (N14493, N14490);
xor XOR2 (N14494, N14486, N4381);
buf BUF1 (N14495, N14478);
nor NOR4 (N14496, N14495, N10177, N3112, N8469);
and AND3 (N14497, N14484, N8721, N8529);
nor NOR3 (N14498, N14487, N6637, N10814);
buf BUF1 (N14499, N14496);
nand NAND2 (N14500, N14485, N14150);
or OR3 (N14501, N14481, N3542, N1764);
buf BUF1 (N14502, N14491);
nor NOR3 (N14503, N14498, N6739, N3674);
nor NOR4 (N14504, N14501, N12188, N8408, N10147);
buf BUF1 (N14505, N14492);
and AND4 (N14506, N14497, N2844, N8098, N7545);
and AND4 (N14507, N14503, N4053, N8367, N8407);
nand NAND3 (N14508, N14493, N13713, N251);
nand NAND2 (N14509, N14506, N14022);
or OR4 (N14510, N14502, N5851, N1559, N6904);
buf BUF1 (N14511, N14499);
xor XOR2 (N14512, N14500, N4004);
not NOT1 (N14513, N14494);
and AND4 (N14514, N14508, N27, N6463, N8287);
and AND4 (N14515, N14511, N4324, N10839, N8833);
and AND3 (N14516, N14509, N42, N14453);
and AND4 (N14517, N14505, N6877, N3493, N7251);
and AND2 (N14518, N14466, N11966);
or OR4 (N14519, N14512, N6496, N10779, N11651);
not NOT1 (N14520, N14519);
and AND4 (N14521, N14520, N10765, N6693, N6202);
and AND3 (N14522, N14510, N6947, N12790);
xor XOR2 (N14523, N14504, N9528);
not NOT1 (N14524, N14521);
xor XOR2 (N14525, N14524, N123);
or OR4 (N14526, N14523, N13892, N13023, N3684);
not NOT1 (N14527, N14518);
or OR3 (N14528, N14517, N9607, N13567);
or OR3 (N14529, N14527, N11047, N10951);
nor NOR4 (N14530, N14522, N7966, N4936, N13767);
nor NOR3 (N14531, N14514, N2725, N14416);
not NOT1 (N14532, N14515);
xor XOR2 (N14533, N14516, N6101);
not NOT1 (N14534, N14526);
and AND3 (N14535, N14531, N4974, N689);
not NOT1 (N14536, N14532);
xor XOR2 (N14537, N14536, N9109);
and AND4 (N14538, N14535, N2195, N6063, N9028);
buf BUF1 (N14539, N14530);
not NOT1 (N14540, N14529);
buf BUF1 (N14541, N14538);
or OR3 (N14542, N14528, N3922, N5016);
nor NOR2 (N14543, N14534, N5239);
not NOT1 (N14544, N14539);
xor XOR2 (N14545, N14533, N11524);
or OR3 (N14546, N14542, N4584, N1895);
or OR3 (N14547, N14544, N3162, N7556);
nand NAND3 (N14548, N14543, N10953, N2965);
nor NOR4 (N14549, N14537, N3690, N8481, N2866);
and AND3 (N14550, N14507, N5468, N10841);
xor XOR2 (N14551, N14547, N13796);
xor XOR2 (N14552, N14540, N5654);
nand NAND3 (N14553, N14513, N9749, N11714);
nand NAND2 (N14554, N14550, N2956);
nor NOR4 (N14555, N14545, N14008, N2698, N224);
not NOT1 (N14556, N14549);
nand NAND3 (N14557, N14541, N487, N6211);
xor XOR2 (N14558, N14556, N10756);
nand NAND2 (N14559, N14558, N5545);
nor NOR3 (N14560, N14557, N8022, N3892);
or OR4 (N14561, N14548, N12612, N2950, N5126);
xor XOR2 (N14562, N14561, N14309);
or OR4 (N14563, N14525, N5826, N14001, N3495);
xor XOR2 (N14564, N14563, N7798);
buf BUF1 (N14565, N14554);
or OR3 (N14566, N14560, N5207, N8146);
buf BUF1 (N14567, N14566);
buf BUF1 (N14568, N14567);
buf BUF1 (N14569, N14555);
and AND2 (N14570, N14565, N4255);
nor NOR3 (N14571, N14559, N8269, N13612);
and AND3 (N14572, N14562, N12383, N12690);
and AND2 (N14573, N14569, N13281);
xor XOR2 (N14574, N14568, N858);
not NOT1 (N14575, N14574);
nand NAND4 (N14576, N14570, N10599, N5485, N11391);
or OR2 (N14577, N14546, N6541);
and AND3 (N14578, N14552, N4883, N7157);
nand NAND3 (N14579, N14572, N6109, N7907);
not NOT1 (N14580, N14575);
or OR4 (N14581, N14553, N11910, N7417, N5844);
buf BUF1 (N14582, N14571);
nand NAND3 (N14583, N14564, N4427, N11633);
nor NOR4 (N14584, N14580, N8242, N1412, N2785);
nor NOR2 (N14585, N14577, N10260);
nand NAND4 (N14586, N14585, N9201, N14540, N203);
not NOT1 (N14587, N14583);
nor NOR4 (N14588, N14582, N13857, N2925, N8941);
nor NOR4 (N14589, N14588, N10270, N1996, N12999);
buf BUF1 (N14590, N14578);
nand NAND2 (N14591, N14579, N4448);
nand NAND4 (N14592, N14573, N10863, N14272, N4022);
xor XOR2 (N14593, N14591, N9187);
or OR4 (N14594, N14581, N10843, N12752, N12298);
or OR4 (N14595, N14576, N10200, N11757, N1871);
or OR4 (N14596, N14593, N8349, N1796, N12140);
nand NAND4 (N14597, N14592, N12667, N10164, N3963);
xor XOR2 (N14598, N14589, N7153);
nor NOR4 (N14599, N14595, N1330, N1921, N2247);
and AND4 (N14600, N14551, N8504, N3187, N13088);
or OR4 (N14601, N14596, N5562, N382, N5539);
nand NAND3 (N14602, N14594, N7393, N12230);
xor XOR2 (N14603, N14601, N9971);
and AND4 (N14604, N14584, N11095, N12394, N2801);
or OR3 (N14605, N14599, N348, N3807);
buf BUF1 (N14606, N14605);
nand NAND3 (N14607, N14600, N10335, N2928);
nand NAND2 (N14608, N14606, N10842);
nor NOR4 (N14609, N14608, N9720, N13454, N10641);
nor NOR3 (N14610, N14609, N8546, N7461);
buf BUF1 (N14611, N14598);
not NOT1 (N14612, N14590);
nor NOR3 (N14613, N14604, N4537, N8807);
or OR3 (N14614, N14610, N1857, N6721);
not NOT1 (N14615, N14607);
xor XOR2 (N14616, N14611, N4214);
nand NAND4 (N14617, N14612, N4040, N10298, N1084);
nand NAND4 (N14618, N14613, N3622, N3906, N4507);
nand NAND4 (N14619, N14614, N1217, N8060, N14421);
and AND2 (N14620, N14616, N12002);
nor NOR4 (N14621, N14602, N8806, N9032, N7283);
buf BUF1 (N14622, N14597);
nand NAND4 (N14623, N14621, N6788, N6023, N13577);
nor NOR4 (N14624, N14587, N5948, N4616, N11410);
not NOT1 (N14625, N14620);
buf BUF1 (N14626, N14615);
buf BUF1 (N14627, N14624);
nand NAND4 (N14628, N14586, N5692, N13771, N7657);
xor XOR2 (N14629, N14603, N8530);
not NOT1 (N14630, N14618);
nand NAND3 (N14631, N14628, N8030, N12976);
nand NAND4 (N14632, N14622, N3173, N11750, N13347);
nor NOR3 (N14633, N14625, N8514, N8639);
nor NOR3 (N14634, N14627, N7130, N4279);
xor XOR2 (N14635, N14617, N14013);
nor NOR3 (N14636, N14631, N11207, N9086);
nor NOR2 (N14637, N14630, N1219);
not NOT1 (N14638, N14636);
nor NOR3 (N14639, N14626, N14047, N7983);
buf BUF1 (N14640, N14635);
xor XOR2 (N14641, N14619, N8688);
or OR3 (N14642, N14632, N9656, N11166);
not NOT1 (N14643, N14637);
buf BUF1 (N14644, N14638);
nand NAND2 (N14645, N14640, N8281);
nand NAND4 (N14646, N14643, N14548, N10928, N6526);
buf BUF1 (N14647, N14644);
nand NAND4 (N14648, N14633, N13573, N2541, N8802);
nor NOR2 (N14649, N14641, N13147);
xor XOR2 (N14650, N14646, N6046);
and AND2 (N14651, N14634, N2267);
or OR4 (N14652, N14629, N3045, N10037, N10098);
nand NAND2 (N14653, N14648, N3854);
and AND2 (N14654, N14650, N6386);
xor XOR2 (N14655, N14651, N7284);
nor NOR2 (N14656, N14642, N8123);
and AND4 (N14657, N14623, N2955, N781, N13982);
or OR4 (N14658, N14639, N8201, N870, N8180);
nor NOR4 (N14659, N14645, N9837, N6969, N1132);
not NOT1 (N14660, N14658);
buf BUF1 (N14661, N14659);
or OR4 (N14662, N14647, N9779, N11572, N2542);
and AND4 (N14663, N14661, N163, N1522, N10690);
xor XOR2 (N14664, N14654, N4871);
and AND2 (N14665, N14649, N12048);
or OR4 (N14666, N14655, N10063, N3952, N8180);
nor NOR2 (N14667, N14653, N7441);
xor XOR2 (N14668, N14667, N5909);
nand NAND4 (N14669, N14656, N13147, N7368, N14533);
nand NAND2 (N14670, N14662, N11085);
not NOT1 (N14671, N14669);
buf BUF1 (N14672, N14670);
xor XOR2 (N14673, N14671, N543);
buf BUF1 (N14674, N14668);
buf BUF1 (N14675, N14663);
not NOT1 (N14676, N14660);
not NOT1 (N14677, N14672);
xor XOR2 (N14678, N14652, N48);
buf BUF1 (N14679, N14678);
xor XOR2 (N14680, N14674, N7428);
nor NOR3 (N14681, N14665, N10826, N3479);
and AND3 (N14682, N14675, N13912, N1437);
xor XOR2 (N14683, N14682, N10114);
nand NAND3 (N14684, N14673, N12985, N10027);
nor NOR3 (N14685, N14666, N4946, N8606);
buf BUF1 (N14686, N14657);
buf BUF1 (N14687, N14677);
nor NOR4 (N14688, N14687, N14662, N9628, N1070);
buf BUF1 (N14689, N14684);
buf BUF1 (N14690, N14664);
xor XOR2 (N14691, N14679, N11406);
nor NOR2 (N14692, N14683, N4414);
xor XOR2 (N14693, N14691, N5744);
and AND3 (N14694, N14681, N5750, N8511);
or OR2 (N14695, N14688, N6741);
xor XOR2 (N14696, N14680, N10323);
or OR2 (N14697, N14695, N9211);
buf BUF1 (N14698, N14696);
nor NOR3 (N14699, N14692, N8585, N7669);
xor XOR2 (N14700, N14694, N10359);
nor NOR2 (N14701, N14699, N9017);
buf BUF1 (N14702, N14701);
or OR3 (N14703, N14690, N14502, N3244);
buf BUF1 (N14704, N14693);
and AND4 (N14705, N14702, N12597, N14377, N14053);
not NOT1 (N14706, N14686);
or OR3 (N14707, N14703, N8082, N7781);
or OR3 (N14708, N14697, N14629, N5276);
xor XOR2 (N14709, N14705, N4764);
buf BUF1 (N14710, N14704);
buf BUF1 (N14711, N14689);
nand NAND3 (N14712, N14676, N7949, N2992);
and AND3 (N14713, N14711, N11326, N12356);
buf BUF1 (N14714, N14708);
nand NAND4 (N14715, N14709, N1006, N2641, N7287);
xor XOR2 (N14716, N14707, N4168);
xor XOR2 (N14717, N14710, N7057);
xor XOR2 (N14718, N14706, N5783);
xor XOR2 (N14719, N14700, N8168);
not NOT1 (N14720, N14716);
buf BUF1 (N14721, N14714);
nand NAND2 (N14722, N14715, N2608);
xor XOR2 (N14723, N14722, N12168);
or OR2 (N14724, N14717, N12504);
buf BUF1 (N14725, N14685);
nand NAND4 (N14726, N14723, N4884, N11445, N10431);
xor XOR2 (N14727, N14719, N13151);
xor XOR2 (N14728, N14712, N1587);
nand NAND3 (N14729, N14727, N13293, N559);
nor NOR4 (N14730, N14728, N9488, N7966, N7315);
nor NOR3 (N14731, N14724, N9953, N9716);
or OR4 (N14732, N14718, N11902, N8989, N8086);
xor XOR2 (N14733, N14732, N8344);
not NOT1 (N14734, N14713);
buf BUF1 (N14735, N14721);
xor XOR2 (N14736, N14720, N4084);
buf BUF1 (N14737, N14731);
buf BUF1 (N14738, N14698);
xor XOR2 (N14739, N14736, N2533);
buf BUF1 (N14740, N14733);
xor XOR2 (N14741, N14725, N7857);
or OR2 (N14742, N14729, N4363);
nor NOR4 (N14743, N14737, N1291, N2590, N13270);
xor XOR2 (N14744, N14735, N6346);
nor NOR4 (N14745, N14742, N1869, N3548, N3226);
not NOT1 (N14746, N14740);
not NOT1 (N14747, N14745);
nor NOR2 (N14748, N14739, N13360);
xor XOR2 (N14749, N14741, N10287);
or OR2 (N14750, N14746, N4618);
buf BUF1 (N14751, N14744);
and AND4 (N14752, N14738, N5874, N1986, N5439);
and AND4 (N14753, N14730, N2139, N2740, N11700);
xor XOR2 (N14754, N14747, N14633);
nand NAND2 (N14755, N14743, N150);
nand NAND3 (N14756, N14749, N12035, N14239);
not NOT1 (N14757, N14752);
xor XOR2 (N14758, N14734, N3626);
xor XOR2 (N14759, N14753, N13299);
buf BUF1 (N14760, N14757);
and AND3 (N14761, N14760, N5143, N6011);
xor XOR2 (N14762, N14761, N8041);
buf BUF1 (N14763, N14754);
and AND3 (N14764, N14726, N13227, N6220);
and AND2 (N14765, N14764, N9886);
buf BUF1 (N14766, N14750);
buf BUF1 (N14767, N14765);
nor NOR2 (N14768, N14751, N134);
and AND4 (N14769, N14759, N10660, N3554, N4679);
or OR2 (N14770, N14768, N12994);
not NOT1 (N14771, N14762);
buf BUF1 (N14772, N14771);
not NOT1 (N14773, N14756);
and AND2 (N14774, N14772, N2169);
xor XOR2 (N14775, N14774, N6486);
xor XOR2 (N14776, N14767, N8713);
nor NOR3 (N14777, N14770, N7464, N8706);
xor XOR2 (N14778, N14758, N11569);
and AND4 (N14779, N14775, N12668, N13107, N3884);
nand NAND2 (N14780, N14778, N14265);
xor XOR2 (N14781, N14763, N8450);
buf BUF1 (N14782, N14780);
not NOT1 (N14783, N14781);
not NOT1 (N14784, N14766);
nor NOR3 (N14785, N14776, N6469, N7665);
not NOT1 (N14786, N14748);
and AND3 (N14787, N14779, N4112, N6890);
not NOT1 (N14788, N14777);
xor XOR2 (N14789, N14787, N10797);
and AND2 (N14790, N14788, N14416);
not NOT1 (N14791, N14782);
not NOT1 (N14792, N14769);
and AND4 (N14793, N14785, N1510, N1041, N4697);
or OR4 (N14794, N14792, N3568, N14508, N9170);
nand NAND2 (N14795, N14790, N6219);
or OR4 (N14796, N14786, N3293, N1811, N6992);
and AND2 (N14797, N14793, N1259);
and AND4 (N14798, N14791, N3686, N8881, N2118);
and AND3 (N14799, N14755, N11356, N1258);
nor NOR3 (N14800, N14798, N9305, N3892);
not NOT1 (N14801, N14797);
nand NAND2 (N14802, N14773, N5542);
nor NOR4 (N14803, N14789, N8080, N10673, N8827);
xor XOR2 (N14804, N14801, N4274);
or OR3 (N14805, N14800, N1498, N14717);
and AND4 (N14806, N14802, N7261, N12882, N13003);
nand NAND2 (N14807, N14794, N182);
xor XOR2 (N14808, N14807, N1449);
xor XOR2 (N14809, N14803, N3743);
or OR4 (N14810, N14809, N13858, N1481, N2247);
or OR3 (N14811, N14810, N7847, N9943);
xor XOR2 (N14812, N14799, N7782);
nand NAND3 (N14813, N14783, N4296, N14591);
and AND3 (N14814, N14811, N8656, N13712);
and AND3 (N14815, N14813, N84, N4496);
buf BUF1 (N14816, N14784);
buf BUF1 (N14817, N14816);
nand NAND4 (N14818, N14805, N6724, N4268, N7291);
buf BUF1 (N14819, N14812);
not NOT1 (N14820, N14806);
nor NOR3 (N14821, N14817, N13173, N7977);
nand NAND3 (N14822, N14796, N142, N9980);
buf BUF1 (N14823, N14819);
or OR4 (N14824, N14804, N13612, N7300, N13414);
or OR3 (N14825, N14818, N9005, N1725);
buf BUF1 (N14826, N14814);
not NOT1 (N14827, N14823);
or OR3 (N14828, N14825, N6340, N9782);
and AND4 (N14829, N14827, N6866, N2540, N10116);
nor NOR3 (N14830, N14808, N12579, N12205);
nor NOR2 (N14831, N14821, N501);
or OR3 (N14832, N14795, N10182, N8848);
xor XOR2 (N14833, N14815, N249);
buf BUF1 (N14834, N14830);
nand NAND2 (N14835, N14832, N4367);
nor NOR2 (N14836, N14829, N3202);
or OR4 (N14837, N14824, N8269, N5609, N3271);
xor XOR2 (N14838, N14826, N5587);
xor XOR2 (N14839, N14834, N4443);
xor XOR2 (N14840, N14828, N9951);
not NOT1 (N14841, N14838);
buf BUF1 (N14842, N14839);
not NOT1 (N14843, N14836);
and AND2 (N14844, N14835, N4074);
buf BUF1 (N14845, N14837);
and AND3 (N14846, N14831, N9381, N10864);
nor NOR2 (N14847, N14844, N3569);
xor XOR2 (N14848, N14847, N3996);
buf BUF1 (N14849, N14848);
xor XOR2 (N14850, N14833, N13117);
or OR4 (N14851, N14820, N5456, N6804, N12063);
nand NAND4 (N14852, N14840, N10777, N14752, N1936);
or OR4 (N14853, N14849, N2089, N5327, N2986);
nor NOR2 (N14854, N14843, N5929);
nor NOR3 (N14855, N14853, N11560, N9119);
not NOT1 (N14856, N14845);
buf BUF1 (N14857, N14854);
not NOT1 (N14858, N14851);
xor XOR2 (N14859, N14822, N12265);
nand NAND2 (N14860, N14856, N727);
nor NOR2 (N14861, N14846, N8402);
buf BUF1 (N14862, N14855);
nor NOR3 (N14863, N14850, N7079, N10310);
buf BUF1 (N14864, N14862);
nand NAND4 (N14865, N14857, N9688, N14803, N8655);
and AND4 (N14866, N14865, N11430, N7333, N3406);
or OR2 (N14867, N14858, N4065);
and AND4 (N14868, N14841, N831, N13098, N9306);
nand NAND3 (N14869, N14852, N2749, N99);
nor NOR4 (N14870, N14859, N7815, N7859, N238);
nor NOR4 (N14871, N14863, N13282, N970, N11464);
nor NOR3 (N14872, N14861, N3302, N3042);
xor XOR2 (N14873, N14866, N2573);
nand NAND4 (N14874, N14871, N13221, N3286, N1847);
buf BUF1 (N14875, N14872);
xor XOR2 (N14876, N14864, N14429);
nor NOR4 (N14877, N14876, N11351, N14760, N1664);
nand NAND4 (N14878, N14842, N10017, N8852, N3976);
not NOT1 (N14879, N14877);
and AND3 (N14880, N14860, N10129, N4693);
buf BUF1 (N14881, N14878);
or OR2 (N14882, N14869, N957);
or OR2 (N14883, N14867, N3021);
buf BUF1 (N14884, N14874);
and AND3 (N14885, N14882, N2190, N14132);
or OR4 (N14886, N14883, N2832, N12395, N2326);
nor NOR4 (N14887, N14881, N1119, N10128, N7646);
not NOT1 (N14888, N14868);
xor XOR2 (N14889, N14885, N11849);
nor NOR3 (N14890, N14884, N5353, N4599);
and AND4 (N14891, N14870, N4404, N13650, N14590);
or OR2 (N14892, N14889, N3548);
nor NOR3 (N14893, N14879, N5385, N9766);
buf BUF1 (N14894, N14892);
nand NAND4 (N14895, N14887, N3880, N1050, N8304);
xor XOR2 (N14896, N14888, N2488);
xor XOR2 (N14897, N14896, N9748);
or OR2 (N14898, N14894, N9527);
or OR4 (N14899, N14875, N3370, N2246, N1434);
not NOT1 (N14900, N14886);
not NOT1 (N14901, N14890);
nor NOR3 (N14902, N14880, N1237, N1595);
not NOT1 (N14903, N14873);
and AND4 (N14904, N14891, N3633, N11539, N6416);
and AND2 (N14905, N14904, N1063);
buf BUF1 (N14906, N14905);
and AND3 (N14907, N14901, N10537, N3985);
and AND2 (N14908, N14898, N9066);
and AND3 (N14909, N14906, N11605, N11316);
xor XOR2 (N14910, N14902, N569);
and AND4 (N14911, N14893, N5891, N239, N16);
nand NAND4 (N14912, N14907, N8300, N12344, N10953);
not NOT1 (N14913, N14899);
xor XOR2 (N14914, N14900, N2134);
or OR2 (N14915, N14909, N11605);
and AND2 (N14916, N14913, N10816);
or OR2 (N14917, N14912, N14904);
nor NOR2 (N14918, N14914, N14330);
nor NOR3 (N14919, N14916, N4808, N1261);
xor XOR2 (N14920, N14908, N1911);
xor XOR2 (N14921, N14919, N3605);
not NOT1 (N14922, N14921);
or OR3 (N14923, N14920, N3434, N1338);
not NOT1 (N14924, N14911);
buf BUF1 (N14925, N14922);
nor NOR4 (N14926, N14897, N745, N6079, N676);
xor XOR2 (N14927, N14924, N6582);
or OR2 (N14928, N14910, N5141);
or OR3 (N14929, N14925, N764, N14800);
and AND4 (N14930, N14928, N7487, N3988, N6157);
not NOT1 (N14931, N14930);
or OR2 (N14932, N14929, N7365);
nand NAND3 (N14933, N14903, N5962, N525);
not NOT1 (N14934, N14915);
or OR2 (N14935, N14923, N468);
buf BUF1 (N14936, N14931);
nand NAND3 (N14937, N14936, N1530, N6541);
and AND4 (N14938, N14917, N4155, N7198, N7657);
or OR2 (N14939, N14926, N9764);
nor NOR3 (N14940, N14927, N14309, N6819);
xor XOR2 (N14941, N14918, N10982);
buf BUF1 (N14942, N14937);
or OR2 (N14943, N14938, N2083);
and AND3 (N14944, N14932, N14502, N5295);
nand NAND3 (N14945, N14933, N725, N9832);
or OR2 (N14946, N14943, N2720);
and AND2 (N14947, N14934, N11224);
nor NOR3 (N14948, N14895, N291, N14463);
nor NOR4 (N14949, N14948, N13111, N3732, N6915);
buf BUF1 (N14950, N14949);
nor NOR2 (N14951, N14947, N7516);
nor NOR2 (N14952, N14946, N13201);
buf BUF1 (N14953, N14939);
nor NOR2 (N14954, N14944, N8503);
or OR2 (N14955, N14950, N76);
or OR3 (N14956, N14954, N8406, N1584);
and AND2 (N14957, N14953, N10887);
nor NOR2 (N14958, N14941, N1826);
not NOT1 (N14959, N14955);
and AND2 (N14960, N14957, N7429);
nor NOR4 (N14961, N14952, N484, N10432, N9852);
xor XOR2 (N14962, N14958, N2690);
nand NAND3 (N14963, N14959, N9677, N14896);
nand NAND4 (N14964, N14945, N11193, N2682, N2629);
nor NOR3 (N14965, N14964, N14009, N9122);
xor XOR2 (N14966, N14962, N9925);
buf BUF1 (N14967, N14961);
or OR4 (N14968, N14967, N3804, N11161, N4140);
xor XOR2 (N14969, N14951, N11211);
buf BUF1 (N14970, N14968);
buf BUF1 (N14971, N14966);
and AND2 (N14972, N14960, N4301);
or OR3 (N14973, N14935, N11172, N9405);
nand NAND2 (N14974, N14956, N3449);
nor NOR3 (N14975, N14971, N13341, N10762);
and AND2 (N14976, N14963, N4186);
nand NAND4 (N14977, N14970, N6174, N8743, N2818);
not NOT1 (N14978, N14969);
nand NAND4 (N14979, N14977, N2496, N9089, N9114);
and AND4 (N14980, N14965, N13874, N14317, N2839);
or OR2 (N14981, N14978, N14298);
or OR4 (N14982, N14973, N11929, N14354, N10529);
buf BUF1 (N14983, N14975);
xor XOR2 (N14984, N14981, N14981);
xor XOR2 (N14985, N14940, N6058);
and AND2 (N14986, N14974, N120);
or OR3 (N14987, N14984, N3603, N8858);
buf BUF1 (N14988, N14979);
xor XOR2 (N14989, N14987, N9529);
and AND3 (N14990, N14983, N9502, N11075);
buf BUF1 (N14991, N14990);
and AND2 (N14992, N14986, N447);
nor NOR3 (N14993, N14985, N12909, N6997);
nand NAND2 (N14994, N14976, N10841);
nand NAND4 (N14995, N14992, N4070, N6204, N6365);
buf BUF1 (N14996, N14982);
buf BUF1 (N14997, N14991);
and AND3 (N14998, N14996, N4938, N316);
xor XOR2 (N14999, N14989, N9269);
not NOT1 (N15000, N14994);
nor NOR3 (N15001, N14942, N10113, N7972);
or OR3 (N15002, N15000, N10444, N8606);
or OR4 (N15003, N14988, N8740, N11894, N4890);
buf BUF1 (N15004, N14993);
buf BUF1 (N15005, N14997);
and AND3 (N15006, N14999, N12215, N1015);
and AND3 (N15007, N15005, N90, N3354);
nand NAND2 (N15008, N15001, N13251);
xor XOR2 (N15009, N14980, N4877);
and AND3 (N15010, N15009, N5809, N11987);
nand NAND4 (N15011, N15003, N10831, N9556, N4630);
and AND3 (N15012, N15011, N5059, N13673);
buf BUF1 (N15013, N15010);
or OR3 (N15014, N15012, N2386, N1495);
and AND2 (N15015, N15014, N1967);
nand NAND2 (N15016, N15004, N11514);
nand NAND4 (N15017, N15007, N9300, N14671, N509);
nor NOR3 (N15018, N15008, N6940, N9047);
nand NAND3 (N15019, N15002, N389, N1163);
xor XOR2 (N15020, N15006, N6399);
and AND3 (N15021, N14972, N12356, N12646);
and AND4 (N15022, N15021, N1772, N2470, N9781);
nor NOR2 (N15023, N15013, N5054);
nand NAND4 (N15024, N15020, N4277, N610, N9559);
nand NAND4 (N15025, N15015, N9717, N1969, N12146);
nor NOR3 (N15026, N15017, N13068, N8440);
buf BUF1 (N15027, N15019);
xor XOR2 (N15028, N15024, N5518);
xor XOR2 (N15029, N14995, N2553);
nor NOR3 (N15030, N15018, N4701, N2573);
nor NOR4 (N15031, N15023, N8372, N9145, N3710);
xor XOR2 (N15032, N15030, N2313);
and AND3 (N15033, N15027, N14659, N8261);
xor XOR2 (N15034, N15029, N3803);
xor XOR2 (N15035, N15028, N7261);
not NOT1 (N15036, N15032);
not NOT1 (N15037, N15036);
or OR4 (N15038, N15022, N9972, N3431, N13885);
not NOT1 (N15039, N15038);
nor NOR4 (N15040, N15033, N12313, N13156, N14177);
xor XOR2 (N15041, N15016, N3878);
nand NAND2 (N15042, N14998, N13975);
or OR3 (N15043, N15039, N2360, N2113);
or OR4 (N15044, N15041, N12425, N666, N9888);
buf BUF1 (N15045, N15037);
buf BUF1 (N15046, N15044);
not NOT1 (N15047, N15025);
buf BUF1 (N15048, N15043);
nor NOR3 (N15049, N15048, N2934, N13371);
nor NOR3 (N15050, N15046, N13507, N346);
not NOT1 (N15051, N15026);
and AND2 (N15052, N15047, N3704);
nand NAND4 (N15053, N15031, N9187, N10135, N6982);
buf BUF1 (N15054, N15050);
not NOT1 (N15055, N15045);
nand NAND4 (N15056, N15055, N6303, N8286, N13049);
not NOT1 (N15057, N15042);
and AND2 (N15058, N15040, N9213);
nor NOR2 (N15059, N15052, N3096);
not NOT1 (N15060, N15059);
nand NAND3 (N15061, N15057, N1764, N12622);
xor XOR2 (N15062, N15053, N7095);
or OR3 (N15063, N15060, N14604, N8302);
not NOT1 (N15064, N15054);
buf BUF1 (N15065, N15034);
nand NAND2 (N15066, N15035, N9296);
buf BUF1 (N15067, N15062);
nand NAND4 (N15068, N15066, N14282, N8643, N6568);
or OR3 (N15069, N15068, N5482, N7891);
nand NAND2 (N15070, N15049, N823);
and AND2 (N15071, N15070, N1583);
or OR4 (N15072, N15069, N9055, N9497, N7608);
and AND2 (N15073, N15072, N1108);
nand NAND4 (N15074, N15067, N3113, N13673, N6678);
xor XOR2 (N15075, N15065, N6091);
xor XOR2 (N15076, N15073, N1517);
nor NOR4 (N15077, N15056, N10746, N2064, N12261);
or OR3 (N15078, N15064, N9715, N11314);
nand NAND3 (N15079, N15075, N7421, N10219);
and AND4 (N15080, N15063, N8332, N13434, N7484);
not NOT1 (N15081, N15061);
nor NOR3 (N15082, N15077, N895, N2546);
nand NAND3 (N15083, N15078, N11127, N1108);
not NOT1 (N15084, N15071);
buf BUF1 (N15085, N15082);
not NOT1 (N15086, N15079);
xor XOR2 (N15087, N15083, N7040);
nor NOR2 (N15088, N15074, N77);
xor XOR2 (N15089, N15085, N431);
nor NOR3 (N15090, N15076, N2310, N8114);
xor XOR2 (N15091, N15058, N3591);
xor XOR2 (N15092, N15091, N7468);
buf BUF1 (N15093, N15087);
nand NAND2 (N15094, N15086, N6001);
buf BUF1 (N15095, N15051);
nor NOR4 (N15096, N15081, N1042, N9424, N11544);
not NOT1 (N15097, N15093);
xor XOR2 (N15098, N15089, N8174);
nor NOR2 (N15099, N15092, N9453);
nand NAND3 (N15100, N15088, N13243, N15047);
nand NAND2 (N15101, N15095, N8042);
or OR2 (N15102, N15084, N6171);
nor NOR4 (N15103, N15090, N3311, N13793, N8140);
nand NAND2 (N15104, N15097, N2458);
nor NOR3 (N15105, N15099, N2670, N978);
not NOT1 (N15106, N15105);
not NOT1 (N15107, N15102);
buf BUF1 (N15108, N15101);
not NOT1 (N15109, N15106);
buf BUF1 (N15110, N15104);
not NOT1 (N15111, N15098);
buf BUF1 (N15112, N15111);
and AND3 (N15113, N15107, N9233, N2844);
nand NAND4 (N15114, N15108, N3488, N11771, N8510);
or OR2 (N15115, N15103, N3732);
xor XOR2 (N15116, N15080, N1942);
nand NAND3 (N15117, N15100, N7903, N11101);
nor NOR4 (N15118, N15114, N6025, N7130, N9230);
nor NOR3 (N15119, N15112, N11379, N7154);
buf BUF1 (N15120, N15115);
buf BUF1 (N15121, N15094);
nor NOR4 (N15122, N15110, N13061, N2475, N13904);
not NOT1 (N15123, N15118);
nor NOR4 (N15124, N15109, N6058, N14401, N10407);
not NOT1 (N15125, N15116);
nand NAND2 (N15126, N15123, N13230);
xor XOR2 (N15127, N15117, N6441);
nor NOR3 (N15128, N15126, N5337, N1652);
not NOT1 (N15129, N15125);
not NOT1 (N15130, N15129);
nor NOR4 (N15131, N15130, N11053, N11234, N2055);
and AND2 (N15132, N15122, N6556);
or OR2 (N15133, N15124, N293);
and AND4 (N15134, N15113, N9328, N12123, N5442);
nor NOR4 (N15135, N15119, N4224, N10587, N6057);
xor XOR2 (N15136, N15131, N2337);
xor XOR2 (N15137, N15134, N4019);
nor NOR2 (N15138, N15096, N3131);
and AND3 (N15139, N15135, N10715, N12053);
not NOT1 (N15140, N15132);
nand NAND4 (N15141, N15137, N9509, N10318, N3636);
nand NAND2 (N15142, N15120, N5563);
not NOT1 (N15143, N15140);
not NOT1 (N15144, N15139);
xor XOR2 (N15145, N15133, N195);
not NOT1 (N15146, N15128);
xor XOR2 (N15147, N15138, N6469);
nand NAND2 (N15148, N15146, N4846);
buf BUF1 (N15149, N15121);
nor NOR2 (N15150, N15142, N4346);
xor XOR2 (N15151, N15150, N14089);
nand NAND4 (N15152, N15127, N4285, N9609, N2368);
nor NOR2 (N15153, N15151, N7966);
xor XOR2 (N15154, N15144, N3881);
and AND2 (N15155, N15154, N2803);
xor XOR2 (N15156, N15153, N11890);
nand NAND2 (N15157, N15136, N10830);
or OR4 (N15158, N15155, N11318, N11633, N11314);
buf BUF1 (N15159, N15152);
or OR4 (N15160, N15147, N1902, N7571, N13074);
not NOT1 (N15161, N15157);
not NOT1 (N15162, N15159);
and AND2 (N15163, N15160, N9354);
xor XOR2 (N15164, N15158, N13350);
nor NOR4 (N15165, N15163, N4691, N5719, N3547);
xor XOR2 (N15166, N15148, N4922);
or OR3 (N15167, N15164, N5150, N1878);
buf BUF1 (N15168, N15167);
xor XOR2 (N15169, N15156, N5380);
buf BUF1 (N15170, N15169);
nand NAND4 (N15171, N15145, N10383, N7774, N2920);
buf BUF1 (N15172, N15165);
and AND2 (N15173, N15171, N1918);
xor XOR2 (N15174, N15172, N2472);
nor NOR2 (N15175, N15170, N1950);
buf BUF1 (N15176, N15166);
buf BUF1 (N15177, N15173);
or OR3 (N15178, N15177, N9892, N1939);
or OR4 (N15179, N15143, N10989, N14157, N11399);
not NOT1 (N15180, N15175);
and AND4 (N15181, N15162, N9618, N5139, N7219);
or OR4 (N15182, N15180, N2189, N24, N2184);
and AND2 (N15183, N15168, N12919);
xor XOR2 (N15184, N15183, N2628);
not NOT1 (N15185, N15176);
xor XOR2 (N15186, N15182, N11225);
buf BUF1 (N15187, N15186);
buf BUF1 (N15188, N15174);
nand NAND4 (N15189, N15184, N4283, N3680, N14644);
nand NAND2 (N15190, N15149, N1650);
or OR2 (N15191, N15179, N6956);
and AND4 (N15192, N15185, N5764, N13202, N5313);
nand NAND4 (N15193, N15191, N10618, N7376, N5631);
nand NAND2 (N15194, N15193, N13375);
and AND3 (N15195, N15189, N6992, N6963);
xor XOR2 (N15196, N15192, N2260);
nor NOR2 (N15197, N15141, N12905);
nor NOR2 (N15198, N15161, N3790);
and AND3 (N15199, N15190, N5725, N10952);
xor XOR2 (N15200, N15197, N9653);
not NOT1 (N15201, N15199);
xor XOR2 (N15202, N15195, N9073);
buf BUF1 (N15203, N15196);
xor XOR2 (N15204, N15201, N12932);
or OR4 (N15205, N15198, N5987, N5998, N13835);
nor NOR3 (N15206, N15204, N1212, N5992);
not NOT1 (N15207, N15181);
nor NOR4 (N15208, N15207, N184, N11975, N266);
and AND3 (N15209, N15188, N7651, N5276);
nor NOR4 (N15210, N15205, N2779, N8136, N7212);
nand NAND4 (N15211, N15194, N14576, N1588, N8520);
buf BUF1 (N15212, N15202);
buf BUF1 (N15213, N15210);
not NOT1 (N15214, N15212);
nand NAND4 (N15215, N15206, N12062, N7641, N1978);
buf BUF1 (N15216, N15203);
or OR2 (N15217, N15208, N1453);
nand NAND4 (N15218, N15215, N9335, N14518, N8490);
not NOT1 (N15219, N15213);
nand NAND3 (N15220, N15209, N11961, N11239);
xor XOR2 (N15221, N15211, N3825);
and AND4 (N15222, N15214, N7956, N8408, N12085);
not NOT1 (N15223, N15222);
nand NAND3 (N15224, N15223, N14245, N6031);
nand NAND4 (N15225, N15217, N11798, N229, N8676);
nor NOR2 (N15226, N15178, N10171);
xor XOR2 (N15227, N15221, N9895);
nor NOR3 (N15228, N15216, N12394, N6587);
not NOT1 (N15229, N15224);
nand NAND4 (N15230, N15228, N9185, N11440, N8974);
not NOT1 (N15231, N15219);
not NOT1 (N15232, N15230);
xor XOR2 (N15233, N15229, N2161);
buf BUF1 (N15234, N15200);
or OR2 (N15235, N15226, N6949);
or OR3 (N15236, N15225, N7839, N11557);
buf BUF1 (N15237, N15227);
nand NAND4 (N15238, N15220, N4860, N8174, N4236);
buf BUF1 (N15239, N15235);
and AND2 (N15240, N15233, N1437);
and AND4 (N15241, N15237, N7592, N9680, N3045);
xor XOR2 (N15242, N15241, N5769);
buf BUF1 (N15243, N15234);
nand NAND4 (N15244, N15187, N10368, N736, N14861);
xor XOR2 (N15245, N15232, N13195);
not NOT1 (N15246, N15240);
nor NOR2 (N15247, N15242, N6810);
not NOT1 (N15248, N15245);
buf BUF1 (N15249, N15239);
not NOT1 (N15250, N15231);
not NOT1 (N15251, N15250);
buf BUF1 (N15252, N15246);
or OR4 (N15253, N15244, N12454, N5705, N4975);
buf BUF1 (N15254, N15249);
nand NAND4 (N15255, N15236, N7267, N2604, N5543);
nor NOR3 (N15256, N15247, N3273, N980);
buf BUF1 (N15257, N15255);
or OR4 (N15258, N15248, N9919, N6725, N6870);
and AND4 (N15259, N15256, N2742, N4847, N5413);
nand NAND2 (N15260, N15218, N7957);
xor XOR2 (N15261, N15253, N7778);
xor XOR2 (N15262, N15254, N12039);
buf BUF1 (N15263, N15257);
and AND2 (N15264, N15251, N6800);
and AND2 (N15265, N15259, N14468);
not NOT1 (N15266, N15258);
or OR3 (N15267, N15238, N1320, N9690);
nor NOR4 (N15268, N15263, N8605, N13572, N8961);
and AND2 (N15269, N15266, N10191);
or OR2 (N15270, N15265, N2407);
and AND4 (N15271, N15260, N2191, N11540, N10430);
and AND2 (N15272, N15262, N2210);
buf BUF1 (N15273, N15261);
buf BUF1 (N15274, N15243);
or OR4 (N15275, N15273, N4051, N7922, N8602);
not NOT1 (N15276, N15269);
or OR4 (N15277, N15274, N12855, N2890, N7729);
nand NAND4 (N15278, N15268, N4920, N10380, N2054);
nor NOR2 (N15279, N15275, N12935);
buf BUF1 (N15280, N15276);
and AND3 (N15281, N15270, N3507, N1507);
buf BUF1 (N15282, N15264);
and AND2 (N15283, N15267, N2351);
not NOT1 (N15284, N15271);
nor NOR3 (N15285, N15252, N5334, N1782);
nor NOR2 (N15286, N15281, N2608);
xor XOR2 (N15287, N15282, N9300);
or OR2 (N15288, N15283, N1555);
buf BUF1 (N15289, N15278);
buf BUF1 (N15290, N15284);
xor XOR2 (N15291, N15289, N10208);
and AND3 (N15292, N15291, N11996, N12233);
or OR2 (N15293, N15292, N13374);
or OR4 (N15294, N15285, N5824, N12074, N720);
and AND2 (N15295, N15280, N8565);
not NOT1 (N15296, N15286);
nand NAND4 (N15297, N15294, N13278, N4216, N9982);
nor NOR2 (N15298, N15290, N11648);
nand NAND4 (N15299, N15287, N14663, N2851, N7315);
not NOT1 (N15300, N15299);
xor XOR2 (N15301, N15300, N2125);
buf BUF1 (N15302, N15297);
not NOT1 (N15303, N15298);
nor NOR2 (N15304, N15295, N3503);
or OR4 (N15305, N15288, N14750, N5315, N83);
not NOT1 (N15306, N15304);
nor NOR2 (N15307, N15279, N5900);
xor XOR2 (N15308, N15277, N14840);
and AND4 (N15309, N15293, N11499, N10845, N2906);
xor XOR2 (N15310, N15296, N12258);
not NOT1 (N15311, N15303);
xor XOR2 (N15312, N15311, N2716);
xor XOR2 (N15313, N15310, N12458);
or OR4 (N15314, N15313, N3591, N11838, N7446);
xor XOR2 (N15315, N15309, N14845);
not NOT1 (N15316, N15314);
nor NOR2 (N15317, N15305, N11911);
not NOT1 (N15318, N15301);
nor NOR3 (N15319, N15308, N11153, N8555);
nand NAND2 (N15320, N15307, N8103);
nor NOR2 (N15321, N15320, N12348);
nor NOR4 (N15322, N15315, N917, N531, N13747);
and AND2 (N15323, N15317, N8839);
xor XOR2 (N15324, N15319, N1594);
buf BUF1 (N15325, N15316);
or OR3 (N15326, N15312, N7658, N2057);
buf BUF1 (N15327, N15321);
buf BUF1 (N15328, N15318);
not NOT1 (N15329, N15326);
nand NAND2 (N15330, N15329, N11392);
buf BUF1 (N15331, N15327);
not NOT1 (N15332, N15322);
nand NAND3 (N15333, N15328, N1015, N1712);
xor XOR2 (N15334, N15325, N2055);
or OR4 (N15335, N15272, N4038, N3332, N2250);
nand NAND4 (N15336, N15335, N9953, N14405, N12568);
nor NOR2 (N15337, N15333, N11771);
nor NOR4 (N15338, N15324, N365, N7791, N2559);
and AND3 (N15339, N15306, N9959, N10);
buf BUF1 (N15340, N15330);
not NOT1 (N15341, N15332);
nor NOR2 (N15342, N15302, N12326);
not NOT1 (N15343, N15336);
nor NOR3 (N15344, N15341, N10511, N4127);
nor NOR3 (N15345, N15331, N1378, N4185);
not NOT1 (N15346, N15344);
or OR3 (N15347, N15323, N1013, N9442);
or OR3 (N15348, N15346, N13115, N3820);
and AND4 (N15349, N15345, N696, N11171, N9671);
nand NAND2 (N15350, N15337, N7317);
buf BUF1 (N15351, N15338);
and AND2 (N15352, N15349, N5484);
not NOT1 (N15353, N15340);
nand NAND2 (N15354, N15350, N2140);
nor NOR4 (N15355, N15334, N8754, N14285, N11594);
buf BUF1 (N15356, N15348);
xor XOR2 (N15357, N15339, N5162);
or OR3 (N15358, N15342, N5690, N8681);
xor XOR2 (N15359, N15343, N3980);
buf BUF1 (N15360, N15357);
or OR4 (N15361, N15360, N1658, N573, N10991);
buf BUF1 (N15362, N15359);
or OR4 (N15363, N15361, N13604, N11050, N8067);
buf BUF1 (N15364, N15351);
nor NOR4 (N15365, N15362, N878, N6177, N2545);
and AND2 (N15366, N15354, N14228);
buf BUF1 (N15367, N15347);
buf BUF1 (N15368, N15366);
and AND3 (N15369, N15367, N2722, N3351);
xor XOR2 (N15370, N15352, N9808);
or OR2 (N15371, N15353, N14329);
nor NOR4 (N15372, N15356, N7902, N2292, N4717);
nor NOR2 (N15373, N15370, N4859);
buf BUF1 (N15374, N15363);
nand NAND3 (N15375, N15368, N15337, N957);
nor NOR3 (N15376, N15374, N287, N3145);
nand NAND4 (N15377, N15369, N12362, N9009, N3052);
nor NOR4 (N15378, N15376, N4818, N8326, N10248);
nor NOR3 (N15379, N15355, N1292, N13638);
nand NAND3 (N15380, N15377, N13457, N5608);
nor NOR4 (N15381, N15375, N2156, N7194, N8177);
nand NAND3 (N15382, N15378, N5672, N10268);
buf BUF1 (N15383, N15364);
xor XOR2 (N15384, N15379, N6904);
not NOT1 (N15385, N15358);
nand NAND3 (N15386, N15371, N8853, N14108);
xor XOR2 (N15387, N15383, N8549);
or OR3 (N15388, N15387, N4900, N2116);
nand NAND4 (N15389, N15372, N8223, N97, N13655);
and AND3 (N15390, N15382, N11977, N1337);
nand NAND2 (N15391, N15389, N3758);
not NOT1 (N15392, N15386);
nor NOR3 (N15393, N15385, N15319, N1237);
buf BUF1 (N15394, N15365);
xor XOR2 (N15395, N15392, N9379);
nand NAND3 (N15396, N15394, N556, N8804);
buf BUF1 (N15397, N15396);
not NOT1 (N15398, N15395);
nand NAND2 (N15399, N15393, N8709);
xor XOR2 (N15400, N15380, N13366);
xor XOR2 (N15401, N15390, N6501);
nand NAND2 (N15402, N15399, N10595);
and AND4 (N15403, N15402, N7625, N7440, N2718);
or OR3 (N15404, N15398, N3146, N5754);
not NOT1 (N15405, N15404);
and AND2 (N15406, N15384, N13783);
nor NOR4 (N15407, N15381, N13260, N6229, N12394);
xor XOR2 (N15408, N15403, N4487);
not NOT1 (N15409, N15391);
xor XOR2 (N15410, N15397, N1972);
and AND2 (N15411, N15405, N3663);
and AND2 (N15412, N15406, N8845);
or OR2 (N15413, N15401, N12796);
nand NAND3 (N15414, N15412, N1375, N12132);
nor NOR3 (N15415, N15413, N12876, N6798);
or OR4 (N15416, N15409, N13628, N12104, N10575);
nor NOR4 (N15417, N15407, N14996, N1057, N14573);
xor XOR2 (N15418, N15373, N5582);
or OR4 (N15419, N15418, N11008, N9861, N7595);
not NOT1 (N15420, N15415);
xor XOR2 (N15421, N15411, N11285);
nand NAND3 (N15422, N15408, N15158, N1608);
nor NOR4 (N15423, N15420, N14783, N11940, N475);
or OR3 (N15424, N15423, N11767, N7849);
and AND2 (N15425, N15388, N3247);
and AND4 (N15426, N15417, N7660, N5841, N11624);
xor XOR2 (N15427, N15410, N3175);
xor XOR2 (N15428, N15400, N7788);
not NOT1 (N15429, N15424);
nor NOR4 (N15430, N15425, N5608, N5583, N11283);
nor NOR3 (N15431, N15427, N12657, N692);
xor XOR2 (N15432, N15426, N15367);
nand NAND2 (N15433, N15429, N3088);
nor NOR3 (N15434, N15414, N2811, N13900);
and AND3 (N15435, N15432, N4567, N2406);
nor NOR3 (N15436, N15428, N4944, N10583);
xor XOR2 (N15437, N15431, N8980);
buf BUF1 (N15438, N15430);
xor XOR2 (N15439, N15438, N6064);
and AND4 (N15440, N15421, N5892, N3347, N11591);
and AND4 (N15441, N15422, N13422, N3216, N10624);
buf BUF1 (N15442, N15419);
nor NOR2 (N15443, N15436, N6906);
nand NAND3 (N15444, N15435, N9924, N8068);
xor XOR2 (N15445, N15443, N14794);
xor XOR2 (N15446, N15440, N7927);
or OR4 (N15447, N15446, N1873, N31, N7030);
nor NOR4 (N15448, N15444, N10614, N11353, N1498);
and AND2 (N15449, N15442, N14296);
nand NAND4 (N15450, N15448, N14415, N5727, N5456);
nor NOR2 (N15451, N15416, N4628);
not NOT1 (N15452, N15433);
nor NOR3 (N15453, N15441, N4962, N3870);
buf BUF1 (N15454, N15451);
xor XOR2 (N15455, N15449, N10705);
and AND2 (N15456, N15454, N11285);
and AND2 (N15457, N15452, N5057);
nor NOR2 (N15458, N15457, N11502);
xor XOR2 (N15459, N15434, N895);
buf BUF1 (N15460, N15456);
not NOT1 (N15461, N15458);
xor XOR2 (N15462, N15459, N4905);
xor XOR2 (N15463, N15453, N6721);
nor NOR3 (N15464, N15450, N13071, N4586);
not NOT1 (N15465, N15460);
xor XOR2 (N15466, N15439, N10489);
nand NAND4 (N15467, N15445, N2297, N14132, N6829);
nand NAND3 (N15468, N15467, N12033, N13046);
and AND4 (N15469, N15447, N11730, N5147, N5800);
buf BUF1 (N15470, N15469);
xor XOR2 (N15471, N15437, N9509);
buf BUF1 (N15472, N15455);
nor NOR3 (N15473, N15465, N12572, N2812);
nand NAND4 (N15474, N15472, N4866, N10452, N2021);
xor XOR2 (N15475, N15473, N4715);
and AND4 (N15476, N15475, N4127, N13916, N14064);
nand NAND4 (N15477, N15461, N5010, N2275, N6924);
buf BUF1 (N15478, N15470);
buf BUF1 (N15479, N15462);
or OR2 (N15480, N15476, N2087);
or OR3 (N15481, N15466, N7945, N13471);
nor NOR4 (N15482, N15479, N13659, N13715, N12460);
or OR3 (N15483, N15474, N12754, N7674);
not NOT1 (N15484, N15464);
or OR4 (N15485, N15477, N9149, N13957, N15035);
nor NOR4 (N15486, N15468, N4021, N3840, N3522);
xor XOR2 (N15487, N15480, N12314);
xor XOR2 (N15488, N15486, N9027);
buf BUF1 (N15489, N15484);
xor XOR2 (N15490, N15483, N6894);
xor XOR2 (N15491, N15490, N2405);
or OR3 (N15492, N15491, N8269, N2937);
not NOT1 (N15493, N15485);
not NOT1 (N15494, N15489);
not NOT1 (N15495, N15488);
xor XOR2 (N15496, N15478, N15290);
xor XOR2 (N15497, N15496, N8994);
nand NAND4 (N15498, N15497, N3418, N5948, N7742);
or OR3 (N15499, N15463, N6270, N5506);
buf BUF1 (N15500, N15471);
buf BUF1 (N15501, N15494);
nand NAND3 (N15502, N15498, N828, N12767);
nor NOR2 (N15503, N15499, N6216);
not NOT1 (N15504, N15503);
or OR4 (N15505, N15504, N433, N5886, N15301);
buf BUF1 (N15506, N15482);
and AND2 (N15507, N15506, N6978);
and AND3 (N15508, N15502, N13822, N12603);
buf BUF1 (N15509, N15508);
nand NAND3 (N15510, N15500, N7950, N12386);
and AND3 (N15511, N15509, N3624, N11688);
not NOT1 (N15512, N15492);
buf BUF1 (N15513, N15507);
and AND3 (N15514, N15495, N1075, N931);
buf BUF1 (N15515, N15513);
not NOT1 (N15516, N15501);
nand NAND4 (N15517, N15493, N2616, N7154, N10073);
xor XOR2 (N15518, N15515, N2583);
or OR4 (N15519, N15516, N15112, N4779, N13874);
and AND4 (N15520, N15481, N12714, N1078, N11950);
and AND4 (N15521, N15487, N2118, N6247, N1519);
buf BUF1 (N15522, N15521);
buf BUF1 (N15523, N15510);
buf BUF1 (N15524, N15519);
nor NOR2 (N15525, N15520, N4692);
not NOT1 (N15526, N15512);
or OR3 (N15527, N15523, N7313, N10861);
nor NOR3 (N15528, N15518, N1733, N397);
xor XOR2 (N15529, N15527, N8889);
nor NOR2 (N15530, N15528, N689);
nor NOR3 (N15531, N15511, N8368, N12980);
xor XOR2 (N15532, N15505, N938);
nand NAND3 (N15533, N15526, N10107, N14069);
buf BUF1 (N15534, N15532);
or OR2 (N15535, N15530, N2439);
not NOT1 (N15536, N15514);
buf BUF1 (N15537, N15531);
or OR2 (N15538, N15537, N5661);
nor NOR4 (N15539, N15517, N7572, N2079, N12930);
nand NAND2 (N15540, N15539, N6393);
buf BUF1 (N15541, N15534);
nor NOR4 (N15542, N15541, N12886, N11443, N3935);
or OR2 (N15543, N15536, N7014);
buf BUF1 (N15544, N15542);
or OR3 (N15545, N15538, N6987, N2377);
not NOT1 (N15546, N15535);
xor XOR2 (N15547, N15529, N5148);
buf BUF1 (N15548, N15543);
or OR3 (N15549, N15533, N9917, N13619);
nand NAND2 (N15550, N15540, N11215);
nand NAND4 (N15551, N15548, N5924, N13148, N1209);
not NOT1 (N15552, N15549);
nor NOR3 (N15553, N15522, N816, N14847);
nor NOR3 (N15554, N15547, N4441, N13465);
or OR4 (N15555, N15525, N9104, N11749, N1571);
and AND2 (N15556, N15524, N4540);
and AND3 (N15557, N15545, N12333, N12999);
nor NOR3 (N15558, N15550, N12344, N11522);
not NOT1 (N15559, N15555);
and AND2 (N15560, N15558, N4491);
nand NAND2 (N15561, N15554, N14774);
and AND3 (N15562, N15546, N7554, N7579);
and AND2 (N15563, N15562, N9269);
not NOT1 (N15564, N15544);
xor XOR2 (N15565, N15561, N7179);
xor XOR2 (N15566, N15557, N7476);
xor XOR2 (N15567, N15552, N6622);
not NOT1 (N15568, N15551);
nand NAND2 (N15569, N15566, N12840);
nand NAND3 (N15570, N15559, N10086, N13347);
nand NAND2 (N15571, N15560, N7743);
xor XOR2 (N15572, N15564, N10020);
not NOT1 (N15573, N15563);
and AND4 (N15574, N15565, N1693, N2619, N10194);
and AND2 (N15575, N15572, N10661);
not NOT1 (N15576, N15568);
nand NAND3 (N15577, N15569, N10901, N13521);
and AND4 (N15578, N15577, N7118, N10127, N6053);
nor NOR3 (N15579, N15574, N1893, N1931);
buf BUF1 (N15580, N15578);
buf BUF1 (N15581, N15570);
and AND3 (N15582, N15573, N6689, N2278);
buf BUF1 (N15583, N15580);
nor NOR3 (N15584, N15556, N2848, N15155);
or OR4 (N15585, N15581, N2067, N903, N1280);
xor XOR2 (N15586, N15584, N9852);
not NOT1 (N15587, N15567);
nor NOR2 (N15588, N15579, N12494);
not NOT1 (N15589, N15587);
nor NOR2 (N15590, N15585, N11312);
nand NAND3 (N15591, N15553, N13297, N8635);
nor NOR2 (N15592, N15588, N11352);
and AND4 (N15593, N15575, N7019, N6204, N11856);
and AND4 (N15594, N15592, N8541, N7551, N2112);
xor XOR2 (N15595, N15583, N850);
buf BUF1 (N15596, N15571);
xor XOR2 (N15597, N15596, N2415);
and AND2 (N15598, N15593, N6510);
or OR3 (N15599, N15595, N3811, N13771);
and AND4 (N15600, N15586, N9471, N716, N4926);
buf BUF1 (N15601, N15599);
and AND4 (N15602, N15576, N7605, N4935, N14062);
nor NOR3 (N15603, N15591, N220, N5545);
not NOT1 (N15604, N15602);
or OR4 (N15605, N15582, N1802, N13043, N13778);
buf BUF1 (N15606, N15590);
nand NAND2 (N15607, N15600, N14242);
nor NOR2 (N15608, N15597, N12365);
xor XOR2 (N15609, N15589, N6250);
nor NOR4 (N15610, N15594, N1053, N13332, N8658);
or OR4 (N15611, N15598, N13810, N7009, N4486);
nor NOR2 (N15612, N15608, N7594);
not NOT1 (N15613, N15603);
buf BUF1 (N15614, N15609);
xor XOR2 (N15615, N15606, N6757);
nor NOR2 (N15616, N15605, N9974);
not NOT1 (N15617, N15604);
buf BUF1 (N15618, N15617);
not NOT1 (N15619, N15615);
xor XOR2 (N15620, N15612, N3030);
and AND4 (N15621, N15613, N6376, N8161, N14347);
nand NAND3 (N15622, N15601, N11730, N12827);
not NOT1 (N15623, N15607);
xor XOR2 (N15624, N15611, N309);
or OR4 (N15625, N15622, N13066, N5669, N8300);
not NOT1 (N15626, N15618);
or OR2 (N15627, N15620, N11960);
xor XOR2 (N15628, N15623, N11298);
and AND4 (N15629, N15627, N9299, N5921, N5525);
not NOT1 (N15630, N15610);
nor NOR2 (N15631, N15626, N7443);
and AND3 (N15632, N15631, N1468, N11237);
and AND4 (N15633, N15630, N4923, N13707, N1423);
not NOT1 (N15634, N15632);
and AND3 (N15635, N15621, N10131, N3472);
and AND4 (N15636, N15614, N7210, N742, N7632);
buf BUF1 (N15637, N15616);
nand NAND4 (N15638, N15634, N9937, N15338, N3244);
buf BUF1 (N15639, N15624);
and AND4 (N15640, N15629, N3238, N9525, N796);
xor XOR2 (N15641, N15636, N4495);
not NOT1 (N15642, N15625);
buf BUF1 (N15643, N15635);
not NOT1 (N15644, N15628);
not NOT1 (N15645, N15641);
or OR2 (N15646, N15619, N48);
and AND3 (N15647, N15642, N7487, N8044);
nor NOR3 (N15648, N15633, N11190, N6140);
not NOT1 (N15649, N15638);
nor NOR2 (N15650, N15649, N12764);
nand NAND4 (N15651, N15648, N12539, N2506, N8927);
not NOT1 (N15652, N15645);
buf BUF1 (N15653, N15651);
nand NAND3 (N15654, N15643, N7858, N5308);
nor NOR3 (N15655, N15654, N6051, N5003);
and AND3 (N15656, N15652, N2908, N3482);
not NOT1 (N15657, N15639);
or OR4 (N15658, N15640, N9557, N7584, N6514);
buf BUF1 (N15659, N15653);
xor XOR2 (N15660, N15659, N11418);
nor NOR3 (N15661, N15646, N6084, N3001);
or OR4 (N15662, N15660, N770, N3204, N11624);
not NOT1 (N15663, N15662);
not NOT1 (N15664, N15663);
nand NAND3 (N15665, N15656, N12142, N15039);
nand NAND3 (N15666, N15665, N14214, N13873);
not NOT1 (N15667, N15657);
and AND2 (N15668, N15647, N10316);
nor NOR4 (N15669, N15661, N7472, N12902, N10512);
and AND4 (N15670, N15668, N2095, N9828, N9114);
nand NAND4 (N15671, N15666, N11727, N531, N12498);
xor XOR2 (N15672, N15637, N11056);
and AND3 (N15673, N15650, N3587, N10124);
or OR2 (N15674, N15669, N3164);
buf BUF1 (N15675, N15667);
or OR2 (N15676, N15658, N153);
or OR3 (N15677, N15674, N14057, N14100);
nand NAND4 (N15678, N15655, N12005, N355, N13841);
not NOT1 (N15679, N15664);
buf BUF1 (N15680, N15676);
nor NOR2 (N15681, N15671, N15524);
xor XOR2 (N15682, N15675, N3027);
nand NAND2 (N15683, N15644, N6884);
buf BUF1 (N15684, N15672);
buf BUF1 (N15685, N15680);
nand NAND3 (N15686, N15685, N3736, N15236);
nor NOR4 (N15687, N15678, N12976, N2008, N968);
or OR4 (N15688, N15679, N2327, N13184, N5986);
nor NOR4 (N15689, N15684, N9126, N691, N13651);
nor NOR2 (N15690, N15689, N10625);
buf BUF1 (N15691, N15690);
nor NOR4 (N15692, N15686, N5297, N9146, N3150);
and AND2 (N15693, N15691, N14650);
nand NAND3 (N15694, N15681, N10479, N832);
and AND4 (N15695, N15673, N7822, N12556, N13177);
nand NAND2 (N15696, N15694, N1605);
nand NAND4 (N15697, N15693, N4801, N11021, N9678);
nor NOR3 (N15698, N15695, N4188, N3398);
or OR4 (N15699, N15682, N7121, N10070, N885);
nand NAND4 (N15700, N15692, N4028, N1503, N4994);
buf BUF1 (N15701, N15698);
or OR3 (N15702, N15670, N13517, N9698);
or OR4 (N15703, N15702, N6135, N10341, N12525);
or OR2 (N15704, N15688, N589);
nor NOR3 (N15705, N15700, N12468, N5977);
or OR2 (N15706, N15687, N15365);
buf BUF1 (N15707, N15704);
buf BUF1 (N15708, N15696);
not NOT1 (N15709, N15705);
nand NAND4 (N15710, N15683, N4478, N4374, N14982);
xor XOR2 (N15711, N15706, N6150);
nor NOR4 (N15712, N15708, N13111, N10429, N8527);
nand NAND4 (N15713, N15699, N342, N3977, N12187);
nor NOR2 (N15714, N15709, N8267);
nand NAND2 (N15715, N15697, N14961);
nor NOR4 (N15716, N15703, N6963, N4954, N664);
xor XOR2 (N15717, N15711, N5449);
and AND2 (N15718, N15677, N4625);
nor NOR4 (N15719, N15714, N14610, N8658, N2100);
or OR3 (N15720, N15717, N1990, N7829);
and AND2 (N15721, N15718, N15390);
xor XOR2 (N15722, N15719, N935);
not NOT1 (N15723, N15712);
not NOT1 (N15724, N15715);
or OR2 (N15725, N15713, N8191);
nor NOR2 (N15726, N15722, N7297);
or OR2 (N15727, N15724, N863);
nand NAND2 (N15728, N15707, N2860);
or OR4 (N15729, N15721, N9250, N3959, N3073);
nand NAND4 (N15730, N15727, N11821, N9250, N5750);
buf BUF1 (N15731, N15726);
xor XOR2 (N15732, N15723, N3752);
or OR3 (N15733, N15720, N14010, N113);
nor NOR2 (N15734, N15710, N614);
nand NAND4 (N15735, N15731, N14832, N5828, N4146);
nand NAND2 (N15736, N15725, N6654);
xor XOR2 (N15737, N15716, N8539);
nand NAND4 (N15738, N15733, N13246, N10543, N12477);
nand NAND3 (N15739, N15730, N3887, N5696);
and AND3 (N15740, N15737, N7009, N9545);
nor NOR4 (N15741, N15732, N15525, N6504, N12506);
xor XOR2 (N15742, N15736, N8797);
xor XOR2 (N15743, N15739, N13118);
nor NOR4 (N15744, N15738, N10913, N13819, N13215);
not NOT1 (N15745, N15701);
nand NAND2 (N15746, N15743, N15698);
nor NOR2 (N15747, N15746, N6195);
xor XOR2 (N15748, N15741, N4330);
nor NOR3 (N15749, N15745, N12302, N10797);
xor XOR2 (N15750, N15747, N8951);
or OR4 (N15751, N15749, N13681, N4940, N5665);
nor NOR4 (N15752, N15748, N15214, N2479, N15713);
and AND4 (N15753, N15728, N554, N11533, N15645);
or OR2 (N15754, N15752, N10058);
buf BUF1 (N15755, N15744);
not NOT1 (N15756, N15740);
xor XOR2 (N15757, N15751, N9254);
and AND4 (N15758, N15735, N12109, N3303, N3956);
nand NAND3 (N15759, N15757, N14730, N10848);
and AND4 (N15760, N15734, N1829, N12113, N12502);
and AND4 (N15761, N15729, N2207, N10506, N10345);
xor XOR2 (N15762, N15758, N4888);
or OR3 (N15763, N15756, N10687, N9960);
xor XOR2 (N15764, N15754, N15439);
xor XOR2 (N15765, N15759, N10449);
buf BUF1 (N15766, N15761);
nor NOR4 (N15767, N15742, N8804, N2537, N11899);
nor NOR2 (N15768, N15763, N6655);
or OR2 (N15769, N15765, N10377);
not NOT1 (N15770, N15768);
or OR3 (N15771, N15760, N804, N13447);
nand NAND2 (N15772, N15771, N13811);
or OR4 (N15773, N15766, N9220, N9918, N2292);
nor NOR3 (N15774, N15770, N9082, N11744);
nor NOR2 (N15775, N15769, N7390);
xor XOR2 (N15776, N15775, N3601);
or OR4 (N15777, N15776, N4712, N4778, N245);
and AND3 (N15778, N15753, N4766, N9128);
nand NAND2 (N15779, N15778, N12389);
xor XOR2 (N15780, N15773, N7723);
not NOT1 (N15781, N15780);
and AND4 (N15782, N15781, N1064, N5895, N3581);
xor XOR2 (N15783, N15779, N8628);
and AND2 (N15784, N15762, N5973);
buf BUF1 (N15785, N15772);
buf BUF1 (N15786, N15777);
xor XOR2 (N15787, N15782, N2145);
nand NAND2 (N15788, N15755, N4290);
or OR4 (N15789, N15785, N614, N1981, N1262);
xor XOR2 (N15790, N15750, N10358);
or OR3 (N15791, N15784, N728, N5297);
nor NOR3 (N15792, N15774, N15148, N2653);
and AND4 (N15793, N15787, N9754, N5924, N13775);
xor XOR2 (N15794, N15764, N2468);
nor NOR4 (N15795, N15792, N13273, N14961, N5214);
xor XOR2 (N15796, N15794, N15716);
and AND4 (N15797, N15790, N7174, N9510, N6411);
and AND2 (N15798, N15797, N9591);
buf BUF1 (N15799, N15783);
nand NAND4 (N15800, N15786, N2991, N418, N10076);
or OR3 (N15801, N15798, N6172, N13780);
and AND2 (N15802, N15796, N9935);
and AND2 (N15803, N15802, N11909);
nand NAND2 (N15804, N15800, N13551);
nor NOR2 (N15805, N15789, N15502);
buf BUF1 (N15806, N15805);
or OR4 (N15807, N15806, N2745, N131, N12134);
not NOT1 (N15808, N15801);
not NOT1 (N15809, N15793);
or OR2 (N15810, N15795, N3434);
or OR2 (N15811, N15799, N13256);
not NOT1 (N15812, N15809);
xor XOR2 (N15813, N15803, N5024);
and AND3 (N15814, N15810, N7299, N9226);
and AND3 (N15815, N15767, N959, N8136);
nand NAND2 (N15816, N15811, N15550);
nand NAND4 (N15817, N15804, N2889, N1565, N15729);
or OR3 (N15818, N15813, N10308, N4138);
buf BUF1 (N15819, N15791);
nand NAND4 (N15820, N15788, N13638, N13996, N12289);
nor NOR3 (N15821, N15814, N6068, N9263);
buf BUF1 (N15822, N15821);
nand NAND2 (N15823, N15808, N8327);
and AND2 (N15824, N15816, N2714);
xor XOR2 (N15825, N15823, N2307);
buf BUF1 (N15826, N15815);
xor XOR2 (N15827, N15826, N4776);
or OR2 (N15828, N15818, N10662);
nor NOR4 (N15829, N15822, N10884, N3465, N2921);
or OR2 (N15830, N15817, N6029);
or OR4 (N15831, N15825, N11236, N11836, N9925);
or OR2 (N15832, N15819, N12806);
or OR3 (N15833, N15820, N6402, N12813);
or OR3 (N15834, N15812, N43, N9695);
nor NOR4 (N15835, N15829, N5138, N14079, N2220);
nand NAND2 (N15836, N15824, N3515);
or OR2 (N15837, N15832, N8977);
xor XOR2 (N15838, N15828, N11643);
xor XOR2 (N15839, N15838, N2296);
not NOT1 (N15840, N15827);
and AND4 (N15841, N15831, N515, N5309, N9270);
or OR3 (N15842, N15836, N3783, N5047);
xor XOR2 (N15843, N15839, N7155);
buf BUF1 (N15844, N15835);
not NOT1 (N15845, N15840);
nor NOR2 (N15846, N15830, N7128);
nor NOR2 (N15847, N15842, N9773);
nand NAND2 (N15848, N15834, N7852);
buf BUF1 (N15849, N15837);
nor NOR2 (N15850, N15847, N8717);
nor NOR3 (N15851, N15850, N2307, N4199);
and AND4 (N15852, N15833, N7825, N12581, N10300);
buf BUF1 (N15853, N15844);
nand NAND4 (N15854, N15848, N9595, N14362, N3003);
nand NAND4 (N15855, N15849, N9181, N5803, N12409);
not NOT1 (N15856, N15855);
xor XOR2 (N15857, N15846, N4285);
nor NOR4 (N15858, N15807, N6482, N10504, N4655);
or OR2 (N15859, N15851, N8174);
or OR3 (N15860, N15843, N7764, N10847);
nor NOR3 (N15861, N15845, N3013, N9243);
buf BUF1 (N15862, N15859);
buf BUF1 (N15863, N15856);
and AND4 (N15864, N15863, N5899, N1959, N752);
nor NOR2 (N15865, N15862, N1273);
buf BUF1 (N15866, N15854);
or OR4 (N15867, N15858, N8172, N8859, N14461);
nand NAND3 (N15868, N15861, N7694, N4666);
nor NOR2 (N15869, N15853, N769);
and AND2 (N15870, N15866, N5658);
and AND3 (N15871, N15870, N12857, N13145);
not NOT1 (N15872, N15860);
not NOT1 (N15873, N15867);
nor NOR2 (N15874, N15873, N8897);
or OR3 (N15875, N15841, N7829, N4674);
or OR4 (N15876, N15871, N9550, N10591, N2278);
and AND2 (N15877, N15876, N5670);
or OR4 (N15878, N15875, N11255, N8998, N9448);
not NOT1 (N15879, N15852);
or OR3 (N15880, N15864, N8184, N5714);
or OR3 (N15881, N15877, N3421, N9602);
not NOT1 (N15882, N15865);
or OR2 (N15883, N15878, N1377);
nand NAND4 (N15884, N15872, N11294, N2761, N743);
nand NAND2 (N15885, N15881, N1982);
or OR2 (N15886, N15868, N4242);
and AND3 (N15887, N15884, N7144, N6686);
nand NAND2 (N15888, N15886, N2459);
buf BUF1 (N15889, N15869);
xor XOR2 (N15890, N15885, N10837);
not NOT1 (N15891, N15874);
nand NAND2 (N15892, N15857, N11155);
xor XOR2 (N15893, N15890, N15229);
or OR2 (N15894, N15879, N10582);
and AND4 (N15895, N15892, N14063, N6523, N3386);
buf BUF1 (N15896, N15894);
nor NOR4 (N15897, N15891, N9108, N7646, N867);
nor NOR2 (N15898, N15882, N11525);
or OR3 (N15899, N15883, N11379, N13231);
not NOT1 (N15900, N15898);
and AND2 (N15901, N15899, N1848);
or OR2 (N15902, N15900, N4430);
xor XOR2 (N15903, N15887, N4146);
not NOT1 (N15904, N15896);
and AND2 (N15905, N15903, N10935);
xor XOR2 (N15906, N15902, N9206);
buf BUF1 (N15907, N15904);
nor NOR4 (N15908, N15907, N14641, N6892, N10878);
nand NAND4 (N15909, N15906, N6660, N3031, N9008);
buf BUF1 (N15910, N15888);
buf BUF1 (N15911, N15880);
buf BUF1 (N15912, N15897);
xor XOR2 (N15913, N15889, N14210);
not NOT1 (N15914, N15912);
buf BUF1 (N15915, N15913);
xor XOR2 (N15916, N15910, N15713);
xor XOR2 (N15917, N15911, N4194);
nand NAND3 (N15918, N15905, N255, N9974);
or OR4 (N15919, N15914, N4922, N7142, N12528);
and AND3 (N15920, N15916, N15127, N6780);
nor NOR2 (N15921, N15917, N81);
and AND4 (N15922, N15920, N5680, N8118, N6781);
not NOT1 (N15923, N15909);
not NOT1 (N15924, N15922);
and AND2 (N15925, N15924, N4575);
not NOT1 (N15926, N15901);
nand NAND3 (N15927, N15926, N7552, N7047);
xor XOR2 (N15928, N15893, N4311);
not NOT1 (N15929, N15919);
and AND2 (N15930, N15925, N4042);
and AND4 (N15931, N15921, N12617, N11645, N1257);
nor NOR4 (N15932, N15918, N12665, N11330, N12868);
nand NAND2 (N15933, N15931, N15459);
or OR2 (N15934, N15930, N2662);
and AND2 (N15935, N15928, N14805);
or OR2 (N15936, N15929, N10064);
or OR3 (N15937, N15936, N14163, N13200);
nand NAND4 (N15938, N15933, N3996, N11550, N7264);
buf BUF1 (N15939, N15927);
or OR2 (N15940, N15934, N13576);
nand NAND3 (N15941, N15915, N748, N11973);
or OR2 (N15942, N15895, N10985);
nand NAND4 (N15943, N15923, N734, N3654, N10889);
not NOT1 (N15944, N15935);
nor NOR3 (N15945, N15944, N2102, N2501);
nor NOR3 (N15946, N15945, N333, N7552);
xor XOR2 (N15947, N15941, N3255);
and AND2 (N15948, N15946, N15872);
nor NOR3 (N15949, N15947, N846, N5929);
not NOT1 (N15950, N15908);
and AND3 (N15951, N15948, N15648, N2466);
nand NAND4 (N15952, N15943, N15628, N6916, N4424);
and AND4 (N15953, N15951, N1499, N6740, N7149);
nand NAND2 (N15954, N15950, N10291);
or OR3 (N15955, N15942, N14376, N8090);
or OR3 (N15956, N15939, N11531, N15163);
nand NAND2 (N15957, N15954, N13057);
not NOT1 (N15958, N15955);
and AND4 (N15959, N15938, N13927, N2671, N12522);
or OR3 (N15960, N15957, N4193, N8588);
or OR3 (N15961, N15940, N14550, N2782);
nor NOR4 (N15962, N15960, N1010, N12183, N130);
and AND2 (N15963, N15958, N9531);
nand NAND2 (N15964, N15959, N3567);
nor NOR3 (N15965, N15952, N9305, N8853);
buf BUF1 (N15966, N15963);
and AND3 (N15967, N15961, N9014, N3910);
nand NAND2 (N15968, N15953, N2471);
buf BUF1 (N15969, N15937);
buf BUF1 (N15970, N15962);
buf BUF1 (N15971, N15964);
nand NAND2 (N15972, N15970, N13287);
buf BUF1 (N15973, N15971);
or OR2 (N15974, N15972, N8530);
or OR3 (N15975, N15974, N8743, N15437);
nor NOR3 (N15976, N15969, N3175, N11539);
or OR2 (N15977, N15949, N8132);
nand NAND4 (N15978, N15975, N7855, N7331, N14529);
nor NOR2 (N15979, N15977, N378);
not NOT1 (N15980, N15966);
nor NOR4 (N15981, N15979, N7863, N15024, N7220);
or OR3 (N15982, N15965, N5611, N12126);
or OR4 (N15983, N15973, N6328, N13110, N15178);
nand NAND3 (N15984, N15980, N12461, N2394);
nor NOR2 (N15985, N15956, N7055);
xor XOR2 (N15986, N15982, N354);
not NOT1 (N15987, N15984);
or OR4 (N15988, N15967, N52, N7227, N3852);
and AND3 (N15989, N15981, N9168, N1867);
buf BUF1 (N15990, N15932);
and AND4 (N15991, N15976, N5456, N2694, N14050);
or OR4 (N15992, N15978, N11245, N13847, N4755);
xor XOR2 (N15993, N15987, N11168);
or OR2 (N15994, N15988, N3639);
buf BUF1 (N15995, N15991);
nand NAND3 (N15996, N15994, N2504, N9635);
xor XOR2 (N15997, N15983, N6981);
nand NAND4 (N15998, N15995, N11463, N13766, N1200);
xor XOR2 (N15999, N15997, N8156);
xor XOR2 (N16000, N15968, N12288);
or OR2 (N16001, N15999, N14837);
or OR3 (N16002, N15998, N5137, N6363);
buf BUF1 (N16003, N15996);
nor NOR3 (N16004, N15990, N1918, N13719);
nand NAND3 (N16005, N15986, N517, N6643);
xor XOR2 (N16006, N16005, N6963);
nor NOR3 (N16007, N16004, N4665, N4125);
or OR2 (N16008, N15992, N8495);
nand NAND2 (N16009, N16008, N3378);
xor XOR2 (N16010, N16002, N122);
buf BUF1 (N16011, N16010);
xor XOR2 (N16012, N16009, N14649);
nor NOR2 (N16013, N16007, N15036);
and AND2 (N16014, N16001, N4470);
or OR2 (N16015, N16012, N780);
nor NOR2 (N16016, N16014, N3460);
xor XOR2 (N16017, N15985, N4631);
not NOT1 (N16018, N15989);
xor XOR2 (N16019, N16016, N7643);
not NOT1 (N16020, N16000);
nand NAND4 (N16021, N16020, N880, N9201, N1305);
nand NAND3 (N16022, N16018, N7144, N5123);
buf BUF1 (N16023, N16006);
endmodule