// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23;

output N3998,N4013,N4018,N4021,N4017,N4007,N4022,N4014,N4016,N4023;

nor NOR4 (N24, N3, N23, N12, N1);
nor NOR4 (N25, N4, N8, N2, N11);
xor XOR2 (N26, N21, N2);
or OR4 (N27, N12, N25, N4, N7);
nand NAND3 (N28, N18, N6, N13);
nand NAND3 (N29, N4, N2, N20);
and AND3 (N30, N18, N26, N17);
and AND3 (N31, N4, N12, N26);
nor NOR4 (N32, N8, N12, N21, N1);
and AND3 (N33, N23, N4, N11);
xor XOR2 (N34, N4, N2);
or OR2 (N35, N18, N7);
or OR3 (N36, N30, N4, N6);
nor NOR2 (N37, N27, N13);
buf BUF1 (N38, N37);
buf BUF1 (N39, N32);
nand NAND3 (N40, N35, N30, N5);
xor XOR2 (N41, N28, N11);
xor XOR2 (N42, N31, N28);
nand NAND2 (N43, N39, N22);
xor XOR2 (N44, N38, N14);
nand NAND2 (N45, N29, N25);
not NOT1 (N46, N41);
and AND4 (N47, N36, N19, N44, N31);
nand NAND3 (N48, N28, N31, N43);
and AND2 (N49, N43, N26);
nor NOR3 (N50, N45, N12, N9);
or OR4 (N51, N48, N11, N22, N41);
xor XOR2 (N52, N40, N16);
nor NOR2 (N53, N42, N29);
and AND4 (N54, N34, N10, N39, N34);
nor NOR2 (N55, N53, N49);
buf BUF1 (N56, N7);
or OR2 (N57, N33, N24);
nor NOR2 (N58, N11, N23);
and AND4 (N59, N52, N22, N35, N38);
xor XOR2 (N60, N59, N1);
or OR4 (N61, N47, N10, N39, N33);
and AND2 (N62, N57, N50);
or OR3 (N63, N58, N15, N55);
nor NOR2 (N64, N53, N37);
or OR2 (N65, N57, N34);
or OR4 (N66, N51, N13, N52, N41);
buf BUF1 (N67, N64);
not NOT1 (N68, N56);
xor XOR2 (N69, N67, N31);
not NOT1 (N70, N60);
nand NAND4 (N71, N54, N54, N62, N19);
buf BUF1 (N72, N30);
buf BUF1 (N73, N46);
nor NOR2 (N74, N68, N10);
xor XOR2 (N75, N71, N73);
nor NOR2 (N76, N3, N2);
nand NAND3 (N77, N74, N72, N11);
nand NAND2 (N78, N11, N61);
or OR4 (N79, N39, N75, N34, N5);
buf BUF1 (N80, N18);
nor NOR2 (N81, N69, N72);
not NOT1 (N82, N63);
nand NAND4 (N83, N79, N61, N17, N12);
nand NAND3 (N84, N83, N36, N49);
buf BUF1 (N85, N80);
xor XOR2 (N86, N81, N19);
and AND3 (N87, N82, N37, N13);
nand NAND4 (N88, N76, N81, N28, N86);
buf BUF1 (N89, N11);
or OR3 (N90, N84, N26, N71);
and AND2 (N91, N90, N72);
or OR2 (N92, N70, N81);
nor NOR2 (N93, N92, N83);
nor NOR3 (N94, N88, N62, N65);
or OR3 (N95, N35, N56, N51);
xor XOR2 (N96, N85, N10);
xor XOR2 (N97, N91, N71);
nor NOR2 (N98, N97, N90);
or OR4 (N99, N98, N47, N52, N98);
and AND4 (N100, N94, N16, N33, N64);
and AND2 (N101, N78, N35);
not NOT1 (N102, N95);
and AND2 (N103, N66, N32);
nor NOR2 (N104, N77, N27);
nand NAND3 (N105, N87, N103, N95);
not NOT1 (N106, N82);
buf BUF1 (N107, N105);
nor NOR2 (N108, N93, N107);
not NOT1 (N109, N73);
buf BUF1 (N110, N96);
nand NAND4 (N111, N106, N48, N22, N66);
or OR3 (N112, N100, N83, N73);
nor NOR2 (N113, N109, N6);
xor XOR2 (N114, N89, N5);
nand NAND4 (N115, N111, N25, N37, N59);
nand NAND2 (N116, N112, N106);
or OR4 (N117, N113, N79, N111, N59);
and AND2 (N118, N102, N17);
or OR2 (N119, N101, N37);
nor NOR4 (N120, N118, N107, N8, N103);
nand NAND3 (N121, N108, N70, N108);
buf BUF1 (N122, N121);
or OR4 (N123, N104, N32, N72, N47);
not NOT1 (N124, N116);
not NOT1 (N125, N124);
nor NOR4 (N126, N125, N74, N48, N61);
xor XOR2 (N127, N123, N15);
or OR2 (N128, N126, N121);
buf BUF1 (N129, N110);
buf BUF1 (N130, N99);
not NOT1 (N131, N114);
not NOT1 (N132, N120);
xor XOR2 (N133, N131, N27);
nand NAND2 (N134, N127, N70);
and AND3 (N135, N129, N59, N34);
and AND4 (N136, N117, N99, N70, N116);
nand NAND4 (N137, N122, N3, N47, N82);
and AND2 (N138, N130, N28);
buf BUF1 (N139, N135);
nor NOR4 (N140, N133, N128, N93, N65);
and AND3 (N141, N119, N25, N75);
nor NOR3 (N142, N30, N128, N125);
buf BUF1 (N143, N134);
buf BUF1 (N144, N143);
and AND4 (N145, N144, N125, N127, N127);
nand NAND3 (N146, N136, N80, N41);
and AND2 (N147, N137, N79);
nand NAND4 (N148, N138, N2, N66, N125);
or OR2 (N149, N148, N104);
buf BUF1 (N150, N149);
nor NOR3 (N151, N146, N47, N60);
xor XOR2 (N152, N147, N93);
xor XOR2 (N153, N132, N130);
or OR4 (N154, N140, N31, N45, N76);
buf BUF1 (N155, N141);
nand NAND4 (N156, N153, N5, N3, N77);
nor NOR2 (N157, N151, N6);
xor XOR2 (N158, N155, N102);
nor NOR4 (N159, N145, N50, N115, N140);
nand NAND2 (N160, N64, N47);
nand NAND4 (N161, N158, N85, N69, N12);
and AND2 (N162, N161, N157);
buf BUF1 (N163, N32);
xor XOR2 (N164, N156, N13);
and AND3 (N165, N152, N62, N51);
nand NAND2 (N166, N163, N92);
nor NOR4 (N167, N150, N133, N61, N30);
xor XOR2 (N168, N164, N91);
nor NOR2 (N169, N142, N161);
or OR2 (N170, N159, N132);
nand NAND2 (N171, N166, N56);
or OR4 (N172, N165, N139, N56, N19);
nor NOR4 (N173, N67, N41, N111, N40);
xor XOR2 (N174, N162, N72);
buf BUF1 (N175, N172);
nor NOR3 (N176, N174, N14, N5);
xor XOR2 (N177, N167, N7);
nor NOR2 (N178, N170, N75);
buf BUF1 (N179, N168);
or OR3 (N180, N177, N114, N160);
nand NAND2 (N181, N170, N110);
and AND2 (N182, N178, N121);
nor NOR4 (N183, N182, N61, N85, N37);
not NOT1 (N184, N175);
buf BUF1 (N185, N169);
and AND4 (N186, N183, N75, N154, N157);
buf BUF1 (N187, N64);
buf BUF1 (N188, N171);
nand NAND3 (N189, N185, N183, N130);
nand NAND4 (N190, N186, N126, N120, N119);
not NOT1 (N191, N184);
buf BUF1 (N192, N176);
buf BUF1 (N193, N189);
nand NAND4 (N194, N190, N138, N183, N19);
buf BUF1 (N195, N180);
xor XOR2 (N196, N192, N40);
not NOT1 (N197, N193);
not NOT1 (N198, N196);
and AND3 (N199, N195, N36, N187);
and AND3 (N200, N5, N191, N150);
nand NAND2 (N201, N108, N26);
nor NOR4 (N202, N194, N31, N11, N139);
nand NAND2 (N203, N179, N135);
nand NAND3 (N204, N200, N74, N111);
nand NAND3 (N205, N173, N5, N30);
nor NOR4 (N206, N204, N92, N110, N44);
buf BUF1 (N207, N199);
and AND4 (N208, N197, N99, N33, N103);
not NOT1 (N209, N198);
nand NAND2 (N210, N205, N44);
not NOT1 (N211, N202);
nand NAND4 (N212, N211, N31, N66, N152);
nor NOR2 (N213, N203, N107);
nor NOR4 (N214, N188, N69, N1, N195);
and AND4 (N215, N214, N123, N158, N203);
nor NOR4 (N216, N206, N157, N128, N205);
or OR2 (N217, N215, N134);
xor XOR2 (N218, N213, N166);
nand NAND4 (N219, N212, N94, N80, N17);
xor XOR2 (N220, N181, N14);
nor NOR2 (N221, N218, N108);
nor NOR2 (N222, N201, N93);
buf BUF1 (N223, N208);
xor XOR2 (N224, N207, N201);
and AND2 (N225, N216, N217);
and AND3 (N226, N187, N141, N100);
buf BUF1 (N227, N210);
or OR2 (N228, N226, N163);
nand NAND4 (N229, N221, N184, N82, N128);
buf BUF1 (N230, N209);
not NOT1 (N231, N219);
xor XOR2 (N232, N227, N16);
or OR4 (N233, N223, N159, N182, N3);
nand NAND3 (N234, N231, N109, N205);
buf BUF1 (N235, N232);
not NOT1 (N236, N228);
xor XOR2 (N237, N234, N158);
not NOT1 (N238, N236);
and AND4 (N239, N235, N11, N189, N110);
and AND3 (N240, N222, N214, N188);
not NOT1 (N241, N220);
xor XOR2 (N242, N241, N216);
buf BUF1 (N243, N230);
nor NOR4 (N244, N224, N192, N178, N197);
and AND3 (N245, N244, N186, N8);
or OR2 (N246, N240, N70);
nand NAND2 (N247, N225, N152);
not NOT1 (N248, N243);
or OR2 (N249, N247, N67);
nand NAND3 (N250, N229, N151, N63);
not NOT1 (N251, N237);
buf BUF1 (N252, N248);
nor NOR3 (N253, N238, N4, N25);
buf BUF1 (N254, N249);
nor NOR2 (N255, N239, N9);
not NOT1 (N256, N253);
or OR2 (N257, N256, N7);
xor XOR2 (N258, N254, N76);
and AND2 (N259, N233, N97);
nand NAND2 (N260, N258, N118);
not NOT1 (N261, N250);
buf BUF1 (N262, N260);
buf BUF1 (N263, N245);
or OR2 (N264, N252, N79);
and AND3 (N265, N255, N247, N91);
not NOT1 (N266, N261);
not NOT1 (N267, N262);
and AND3 (N268, N267, N209, N54);
nand NAND3 (N269, N242, N250, N263);
buf BUF1 (N270, N212);
nor NOR3 (N271, N259, N168, N18);
not NOT1 (N272, N246);
or OR3 (N273, N268, N60, N191);
nor NOR4 (N274, N272, N59, N228, N209);
and AND4 (N275, N273, N124, N86, N247);
or OR3 (N276, N270, N275, N14);
and AND2 (N277, N75, N165);
or OR4 (N278, N265, N181, N11, N38);
nand NAND4 (N279, N271, N274, N122, N258);
xor XOR2 (N280, N263, N157);
or OR2 (N281, N251, N223);
nor NOR3 (N282, N280, N189, N137);
nor NOR4 (N283, N279, N177, N264, N261);
not NOT1 (N284, N93);
or OR4 (N285, N283, N127, N12, N76);
not NOT1 (N286, N266);
not NOT1 (N287, N281);
or OR2 (N288, N284, N148);
buf BUF1 (N289, N285);
buf BUF1 (N290, N286);
buf BUF1 (N291, N288);
xor XOR2 (N292, N282, N236);
xor XOR2 (N293, N269, N38);
and AND3 (N294, N290, N158, N243);
xor XOR2 (N295, N291, N272);
xor XOR2 (N296, N276, N3);
nor NOR2 (N297, N287, N48);
xor XOR2 (N298, N295, N112);
nor NOR4 (N299, N296, N83, N294, N280);
and AND3 (N300, N222, N168, N4);
buf BUF1 (N301, N300);
nor NOR4 (N302, N289, N173, N253, N53);
buf BUF1 (N303, N277);
not NOT1 (N304, N298);
not NOT1 (N305, N303);
and AND3 (N306, N293, N146, N108);
nor NOR4 (N307, N305, N35, N99, N290);
buf BUF1 (N308, N299);
xor XOR2 (N309, N308, N252);
and AND2 (N310, N292, N283);
or OR3 (N311, N310, N299, N45);
and AND2 (N312, N301, N299);
not NOT1 (N313, N304);
not NOT1 (N314, N297);
buf BUF1 (N315, N302);
nand NAND4 (N316, N257, N53, N174, N60);
buf BUF1 (N317, N306);
nand NAND4 (N318, N278, N170, N147, N105);
and AND2 (N319, N312, N111);
nor NOR4 (N320, N319, N110, N21, N112);
and AND4 (N321, N314, N225, N107, N23);
nor NOR2 (N322, N309, N184);
or OR3 (N323, N315, N236, N153);
and AND2 (N324, N322, N236);
not NOT1 (N325, N316);
nand NAND4 (N326, N324, N8, N191, N19);
not NOT1 (N327, N311);
not NOT1 (N328, N326);
nand NAND2 (N329, N328, N178);
not NOT1 (N330, N325);
and AND4 (N331, N318, N179, N37, N186);
and AND3 (N332, N329, N308, N271);
buf BUF1 (N333, N321);
nand NAND4 (N334, N313, N153, N123, N10);
nor NOR2 (N335, N330, N188);
nor NOR2 (N336, N320, N173);
xor XOR2 (N337, N331, N248);
buf BUF1 (N338, N333);
xor XOR2 (N339, N327, N222);
nand NAND3 (N340, N317, N249, N246);
nand NAND4 (N341, N340, N191, N70, N116);
or OR4 (N342, N339, N238, N307, N176);
buf BUF1 (N343, N166);
not NOT1 (N344, N323);
or OR2 (N345, N332, N90);
xor XOR2 (N346, N337, N90);
xor XOR2 (N347, N336, N252);
nor NOR2 (N348, N345, N36);
and AND2 (N349, N341, N182);
not NOT1 (N350, N347);
and AND2 (N351, N342, N130);
nand NAND3 (N352, N351, N66, N220);
nor NOR4 (N353, N350, N197, N65, N119);
or OR4 (N354, N352, N131, N353, N321);
nand NAND2 (N355, N111, N109);
and AND2 (N356, N355, N176);
xor XOR2 (N357, N343, N304);
nand NAND2 (N358, N348, N130);
xor XOR2 (N359, N354, N79);
or OR2 (N360, N359, N343);
buf BUF1 (N361, N344);
or OR2 (N362, N349, N190);
not NOT1 (N363, N338);
nand NAND2 (N364, N356, N119);
not NOT1 (N365, N346);
or OR4 (N366, N365, N174, N122, N63);
and AND4 (N367, N362, N62, N265, N222);
nand NAND3 (N368, N357, N44, N141);
nor NOR4 (N369, N366, N318, N207, N329);
buf BUF1 (N370, N358);
and AND3 (N371, N361, N292, N16);
nor NOR2 (N372, N335, N173);
and AND4 (N373, N360, N242, N34, N36);
not NOT1 (N374, N334);
not NOT1 (N375, N364);
and AND3 (N376, N372, N103, N87);
and AND4 (N377, N373, N261, N19, N96);
or OR2 (N378, N370, N303);
nand NAND2 (N379, N367, N283);
nor NOR2 (N380, N369, N134);
xor XOR2 (N381, N376, N288);
xor XOR2 (N382, N375, N307);
nor NOR2 (N383, N374, N331);
nor NOR2 (N384, N383, N51);
not NOT1 (N385, N377);
buf BUF1 (N386, N371);
nand NAND3 (N387, N379, N228, N90);
buf BUF1 (N388, N363);
and AND4 (N389, N378, N101, N67, N19);
and AND2 (N390, N368, N117);
xor XOR2 (N391, N380, N89);
buf BUF1 (N392, N387);
or OR2 (N393, N390, N83);
xor XOR2 (N394, N388, N232);
or OR4 (N395, N382, N64, N387, N192);
and AND2 (N396, N392, N147);
xor XOR2 (N397, N394, N317);
xor XOR2 (N398, N389, N393);
or OR4 (N399, N241, N348, N48, N32);
nor NOR4 (N400, N384, N251, N396, N136);
and AND2 (N401, N321, N300);
not NOT1 (N402, N400);
buf BUF1 (N403, N402);
xor XOR2 (N404, N386, N125);
or OR4 (N405, N401, N117, N204, N145);
not NOT1 (N406, N385);
and AND4 (N407, N403, N402, N348, N361);
nor NOR2 (N408, N391, N84);
buf BUF1 (N409, N395);
buf BUF1 (N410, N404);
buf BUF1 (N411, N399);
buf BUF1 (N412, N381);
not NOT1 (N413, N409);
nor NOR3 (N414, N410, N394, N362);
or OR2 (N415, N412, N318);
nand NAND2 (N416, N408, N19);
and AND3 (N417, N398, N28, N224);
not NOT1 (N418, N397);
nand NAND2 (N419, N415, N172);
xor XOR2 (N420, N416, N94);
buf BUF1 (N421, N414);
and AND3 (N422, N420, N1, N177);
nor NOR3 (N423, N407, N314, N310);
and AND4 (N424, N411, N23, N100, N353);
not NOT1 (N425, N417);
and AND3 (N426, N422, N231, N154);
buf BUF1 (N427, N418);
or OR2 (N428, N426, N162);
nor NOR2 (N429, N425, N221);
nor NOR3 (N430, N427, N57, N317);
nand NAND4 (N431, N406, N284, N367, N384);
and AND3 (N432, N428, N153, N21);
not NOT1 (N433, N423);
not NOT1 (N434, N419);
not NOT1 (N435, N433);
and AND2 (N436, N424, N351);
nor NOR3 (N437, N432, N320, N337);
nor NOR3 (N438, N434, N344, N214);
xor XOR2 (N439, N437, N136);
nand NAND2 (N440, N435, N289);
nand NAND4 (N441, N439, N104, N32, N349);
xor XOR2 (N442, N405, N364);
not NOT1 (N443, N413);
or OR3 (N444, N431, N274, N419);
not NOT1 (N445, N442);
and AND4 (N446, N445, N31, N97, N133);
nand NAND2 (N447, N444, N115);
or OR3 (N448, N447, N90, N191);
not NOT1 (N449, N446);
and AND2 (N450, N438, N145);
nand NAND3 (N451, N440, N378, N124);
xor XOR2 (N452, N451, N80);
nand NAND3 (N453, N429, N266, N144);
buf BUF1 (N454, N441);
not NOT1 (N455, N452);
nand NAND2 (N456, N436, N89);
xor XOR2 (N457, N448, N2);
or OR4 (N458, N456, N380, N292, N92);
and AND4 (N459, N449, N197, N244, N281);
nand NAND4 (N460, N443, N64, N266, N231);
xor XOR2 (N461, N459, N280);
nor NOR3 (N462, N461, N308, N233);
nand NAND4 (N463, N450, N67, N131, N147);
xor XOR2 (N464, N457, N117);
and AND3 (N465, N463, N28, N100);
nand NAND4 (N466, N465, N440, N463, N232);
nor NOR3 (N467, N455, N453, N359);
and AND2 (N468, N333, N96);
not NOT1 (N469, N466);
nand NAND3 (N470, N460, N71, N454);
nor NOR4 (N471, N82, N404, N65, N227);
xor XOR2 (N472, N468, N40);
nor NOR4 (N473, N469, N126, N38, N202);
not NOT1 (N474, N467);
nor NOR2 (N475, N471, N304);
xor XOR2 (N476, N421, N414);
xor XOR2 (N477, N458, N382);
nor NOR2 (N478, N475, N83);
not NOT1 (N479, N474);
not NOT1 (N480, N470);
not NOT1 (N481, N478);
xor XOR2 (N482, N477, N133);
xor XOR2 (N483, N476, N71);
nor NOR4 (N484, N482, N36, N458, N176);
and AND4 (N485, N473, N375, N423, N154);
or OR2 (N486, N464, N413);
or OR2 (N487, N479, N175);
buf BUF1 (N488, N430);
or OR2 (N489, N462, N458);
xor XOR2 (N490, N472, N364);
buf BUF1 (N491, N490);
buf BUF1 (N492, N481);
buf BUF1 (N493, N487);
buf BUF1 (N494, N489);
nand NAND3 (N495, N494, N274, N81);
nor NOR2 (N496, N495, N243);
nand NAND3 (N497, N480, N227, N109);
nand NAND3 (N498, N497, N126, N80);
xor XOR2 (N499, N498, N415);
nand NAND2 (N500, N499, N472);
buf BUF1 (N501, N484);
nand NAND2 (N502, N486, N401);
and AND4 (N503, N491, N243, N280, N240);
buf BUF1 (N504, N500);
or OR4 (N505, N488, N114, N306, N62);
xor XOR2 (N506, N501, N189);
and AND4 (N507, N506, N138, N255, N328);
and AND3 (N508, N483, N458, N87);
buf BUF1 (N509, N485);
nand NAND2 (N510, N507, N96);
not NOT1 (N511, N502);
and AND3 (N512, N504, N224, N86);
xor XOR2 (N513, N512, N373);
and AND2 (N514, N493, N264);
and AND2 (N515, N505, N323);
buf BUF1 (N516, N508);
and AND4 (N517, N510, N263, N462, N439);
xor XOR2 (N518, N509, N378);
nor NOR2 (N519, N513, N207);
xor XOR2 (N520, N496, N71);
and AND4 (N521, N517, N244, N458, N382);
nor NOR2 (N522, N492, N168);
nor NOR4 (N523, N522, N369, N244, N331);
or OR4 (N524, N519, N173, N225, N313);
not NOT1 (N525, N523);
or OR4 (N526, N518, N83, N333, N98);
xor XOR2 (N527, N516, N53);
nand NAND2 (N528, N520, N214);
nand NAND2 (N529, N527, N274);
or OR3 (N530, N503, N148, N451);
nand NAND3 (N531, N529, N358, N297);
or OR4 (N532, N531, N159, N273, N409);
nand NAND2 (N533, N521, N404);
xor XOR2 (N534, N526, N178);
nand NAND2 (N535, N511, N265);
or OR4 (N536, N532, N225, N176, N329);
not NOT1 (N537, N528);
and AND4 (N538, N535, N448, N202, N457);
and AND2 (N539, N514, N239);
xor XOR2 (N540, N534, N251);
xor XOR2 (N541, N538, N432);
and AND3 (N542, N536, N416, N157);
and AND3 (N543, N524, N88, N23);
nor NOR2 (N544, N537, N275);
nand NAND2 (N545, N540, N117);
or OR2 (N546, N545, N233);
xor XOR2 (N547, N530, N43);
or OR3 (N548, N547, N356, N180);
nand NAND3 (N549, N546, N259, N522);
not NOT1 (N550, N548);
nand NAND2 (N551, N525, N167);
nor NOR2 (N552, N515, N25);
or OR3 (N553, N552, N146, N110);
buf BUF1 (N554, N539);
nor NOR3 (N555, N533, N443, N27);
nor NOR2 (N556, N550, N372);
nor NOR2 (N557, N541, N349);
xor XOR2 (N558, N543, N226);
buf BUF1 (N559, N557);
xor XOR2 (N560, N544, N217);
or OR4 (N561, N553, N372, N75, N7);
nand NAND4 (N562, N554, N548, N87, N245);
xor XOR2 (N563, N558, N85);
not NOT1 (N564, N561);
buf BUF1 (N565, N542);
or OR4 (N566, N562, N454, N422, N206);
nor NOR2 (N567, N566, N419);
buf BUF1 (N568, N563);
nand NAND4 (N569, N559, N48, N83, N34);
not NOT1 (N570, N556);
nand NAND3 (N571, N570, N19, N364);
nand NAND2 (N572, N569, N140);
not NOT1 (N573, N560);
nor NOR4 (N574, N568, N28, N192, N490);
and AND2 (N575, N564, N126);
or OR3 (N576, N549, N58, N340);
and AND2 (N577, N572, N179);
or OR3 (N578, N577, N114, N192);
or OR4 (N579, N551, N246, N429, N119);
or OR3 (N580, N579, N421, N26);
or OR4 (N581, N565, N20, N237, N181);
not NOT1 (N582, N555);
or OR4 (N583, N574, N127, N563, N410);
nor NOR2 (N584, N571, N537);
xor XOR2 (N585, N573, N185);
or OR4 (N586, N582, N426, N271, N498);
xor XOR2 (N587, N581, N9);
nor NOR3 (N588, N585, N38, N314);
or OR2 (N589, N578, N489);
or OR2 (N590, N588, N135);
nor NOR4 (N591, N586, N443, N431, N211);
and AND3 (N592, N590, N325, N573);
buf BUF1 (N593, N583);
or OR4 (N594, N593, N112, N41, N18);
or OR2 (N595, N594, N66);
not NOT1 (N596, N567);
nor NOR3 (N597, N592, N546, N38);
or OR4 (N598, N575, N171, N186, N562);
buf BUF1 (N599, N595);
nand NAND4 (N600, N580, N385, N230, N238);
or OR2 (N601, N600, N542);
not NOT1 (N602, N587);
buf BUF1 (N603, N602);
or OR3 (N604, N589, N488, N69);
or OR4 (N605, N584, N72, N330, N530);
buf BUF1 (N606, N597);
buf BUF1 (N607, N599);
and AND2 (N608, N605, N515);
xor XOR2 (N609, N596, N81);
and AND3 (N610, N608, N397, N306);
xor XOR2 (N611, N604, N338);
and AND4 (N612, N610, N581, N371, N495);
nand NAND3 (N613, N598, N379, N409);
buf BUF1 (N614, N607);
xor XOR2 (N615, N576, N520);
nand NAND2 (N616, N606, N76);
nand NAND2 (N617, N616, N381);
not NOT1 (N618, N613);
xor XOR2 (N619, N603, N474);
xor XOR2 (N620, N619, N451);
not NOT1 (N621, N615);
not NOT1 (N622, N601);
nand NAND2 (N623, N591, N277);
or OR3 (N624, N612, N97, N414);
or OR2 (N625, N623, N621);
or OR3 (N626, N176, N374, N385);
nand NAND3 (N627, N611, N218, N557);
and AND2 (N628, N622, N608);
nor NOR2 (N629, N624, N417);
or OR3 (N630, N628, N550, N512);
nor NOR3 (N631, N609, N483, N122);
nand NAND4 (N632, N618, N434, N625, N550);
nand NAND4 (N633, N544, N28, N568, N29);
xor XOR2 (N634, N627, N81);
xor XOR2 (N635, N632, N274);
and AND3 (N636, N630, N274, N569);
xor XOR2 (N637, N634, N469);
and AND4 (N638, N620, N107, N361, N182);
nand NAND4 (N639, N637, N202, N133, N398);
buf BUF1 (N640, N614);
or OR3 (N641, N635, N500, N18);
and AND3 (N642, N639, N166, N574);
not NOT1 (N643, N641);
nand NAND2 (N644, N643, N382);
nor NOR3 (N645, N636, N486, N520);
buf BUF1 (N646, N640);
not NOT1 (N647, N631);
xor XOR2 (N648, N617, N69);
not NOT1 (N649, N642);
nand NAND3 (N650, N629, N461, N533);
nor NOR3 (N651, N626, N383, N527);
xor XOR2 (N652, N644, N122);
xor XOR2 (N653, N645, N382);
nand NAND4 (N654, N646, N84, N262, N235);
buf BUF1 (N655, N633);
buf BUF1 (N656, N652);
and AND2 (N657, N654, N207);
and AND3 (N658, N650, N383, N304);
nor NOR2 (N659, N653, N278);
or OR4 (N660, N655, N397, N87, N418);
not NOT1 (N661, N660);
or OR4 (N662, N638, N602, N348, N187);
xor XOR2 (N663, N651, N303);
nand NAND4 (N664, N647, N325, N225, N498);
not NOT1 (N665, N663);
nand NAND3 (N666, N649, N302, N567);
nand NAND2 (N667, N664, N427);
and AND3 (N668, N667, N120, N45);
or OR4 (N669, N648, N335, N53, N192);
xor XOR2 (N670, N666, N232);
nand NAND3 (N671, N665, N639, N241);
nor NOR3 (N672, N658, N347, N26);
xor XOR2 (N673, N661, N75);
nor NOR2 (N674, N659, N62);
and AND4 (N675, N670, N237, N92, N89);
and AND2 (N676, N674, N253);
not NOT1 (N677, N668);
not NOT1 (N678, N677);
buf BUF1 (N679, N676);
and AND3 (N680, N657, N454, N225);
and AND4 (N681, N673, N294, N288, N186);
not NOT1 (N682, N672);
and AND3 (N683, N678, N280, N60);
xor XOR2 (N684, N683, N132);
and AND2 (N685, N682, N621);
buf BUF1 (N686, N679);
and AND3 (N687, N671, N453, N99);
nand NAND2 (N688, N685, N363);
or OR4 (N689, N688, N191, N425, N646);
buf BUF1 (N690, N662);
nor NOR3 (N691, N690, N622, N468);
nor NOR4 (N692, N669, N639, N435, N452);
xor XOR2 (N693, N686, N98);
xor XOR2 (N694, N681, N82);
or OR2 (N695, N656, N474);
and AND2 (N696, N689, N374);
xor XOR2 (N697, N694, N537);
nor NOR2 (N698, N696, N371);
xor XOR2 (N699, N691, N531);
buf BUF1 (N700, N687);
nand NAND2 (N701, N697, N384);
buf BUF1 (N702, N680);
xor XOR2 (N703, N695, N440);
buf BUF1 (N704, N703);
and AND2 (N705, N701, N596);
nand NAND2 (N706, N705, N344);
buf BUF1 (N707, N693);
and AND2 (N708, N692, N108);
nor NOR4 (N709, N698, N432, N654, N405);
buf BUF1 (N710, N706);
nor NOR3 (N711, N704, N508, N174);
or OR3 (N712, N710, N638, N529);
or OR2 (N713, N702, N292);
and AND2 (N714, N707, N51);
nand NAND2 (N715, N684, N120);
or OR4 (N716, N708, N539, N301, N216);
xor XOR2 (N717, N700, N83);
not NOT1 (N718, N712);
buf BUF1 (N719, N715);
or OR2 (N720, N675, N100);
buf BUF1 (N721, N719);
and AND2 (N722, N717, N691);
or OR3 (N723, N721, N594, N485);
nand NAND4 (N724, N722, N472, N333, N62);
and AND4 (N725, N711, N113, N154, N121);
or OR3 (N726, N709, N105, N238);
nand NAND2 (N727, N720, N258);
and AND2 (N728, N699, N285);
buf BUF1 (N729, N727);
buf BUF1 (N730, N724);
and AND3 (N731, N730, N387, N577);
not NOT1 (N732, N718);
buf BUF1 (N733, N731);
buf BUF1 (N734, N729);
nor NOR3 (N735, N723, N368, N260);
buf BUF1 (N736, N725);
xor XOR2 (N737, N735, N565);
and AND3 (N738, N732, N326, N48);
nand NAND3 (N739, N726, N404, N65);
nor NOR3 (N740, N713, N548, N154);
xor XOR2 (N741, N740, N181);
xor XOR2 (N742, N741, N59);
not NOT1 (N743, N734);
and AND2 (N744, N714, N152);
buf BUF1 (N745, N743);
and AND2 (N746, N728, N105);
and AND4 (N747, N739, N386, N652, N428);
nand NAND4 (N748, N746, N33, N452, N102);
xor XOR2 (N749, N733, N691);
xor XOR2 (N750, N749, N177);
nor NOR3 (N751, N737, N199, N645);
buf BUF1 (N752, N747);
nand NAND4 (N753, N752, N600, N43, N669);
nand NAND3 (N754, N742, N187, N383);
buf BUF1 (N755, N744);
xor XOR2 (N756, N751, N485);
not NOT1 (N757, N756);
xor XOR2 (N758, N716, N33);
xor XOR2 (N759, N750, N304);
not NOT1 (N760, N745);
and AND4 (N761, N760, N673, N603, N735);
buf BUF1 (N762, N754);
nor NOR4 (N763, N762, N739, N669, N402);
nor NOR3 (N764, N748, N73, N423);
buf BUF1 (N765, N758);
or OR3 (N766, N738, N121, N101);
nor NOR2 (N767, N764, N700);
nand NAND2 (N768, N767, N513);
nand NAND3 (N769, N759, N426, N151);
nor NOR3 (N770, N761, N239, N56);
nand NAND2 (N771, N736, N22);
or OR2 (N772, N768, N580);
buf BUF1 (N773, N770);
xor XOR2 (N774, N769, N591);
nand NAND2 (N775, N771, N436);
xor XOR2 (N776, N773, N206);
not NOT1 (N777, N775);
nand NAND2 (N778, N757, N457);
and AND4 (N779, N778, N175, N528, N692);
or OR3 (N780, N763, N229, N299);
buf BUF1 (N781, N753);
or OR4 (N782, N781, N765, N128, N690);
nand NAND2 (N783, N444, N139);
or OR3 (N784, N766, N740, N437);
or OR2 (N785, N777, N427);
nand NAND3 (N786, N784, N566, N366);
or OR2 (N787, N755, N578);
nor NOR2 (N788, N785, N126);
not NOT1 (N789, N772);
buf BUF1 (N790, N787);
and AND2 (N791, N783, N85);
and AND3 (N792, N788, N281, N124);
nand NAND4 (N793, N791, N569, N699, N228);
and AND3 (N794, N776, N235, N549);
nand NAND2 (N795, N790, N719);
xor XOR2 (N796, N786, N507);
and AND3 (N797, N789, N258, N548);
buf BUF1 (N798, N782);
or OR2 (N799, N798, N429);
and AND2 (N800, N794, N648);
nor NOR4 (N801, N779, N353, N262, N784);
or OR3 (N802, N800, N777, N490);
buf BUF1 (N803, N793);
and AND4 (N804, N799, N398, N735, N134);
nor NOR4 (N805, N801, N55, N553, N92);
buf BUF1 (N806, N797);
and AND4 (N807, N774, N654, N276, N92);
buf BUF1 (N808, N796);
not NOT1 (N809, N795);
nor NOR3 (N810, N805, N207, N250);
and AND3 (N811, N803, N314, N180);
xor XOR2 (N812, N811, N89);
not NOT1 (N813, N802);
not NOT1 (N814, N808);
xor XOR2 (N815, N806, N619);
not NOT1 (N816, N792);
nor NOR2 (N817, N804, N697);
nand NAND4 (N818, N812, N283, N810, N373);
and AND3 (N819, N614, N37, N789);
and AND4 (N820, N816, N735, N742, N81);
or OR4 (N821, N814, N170, N122, N36);
nor NOR2 (N822, N821, N114);
nand NAND2 (N823, N818, N422);
not NOT1 (N824, N822);
xor XOR2 (N825, N813, N423);
or OR4 (N826, N824, N345, N571, N273);
nor NOR4 (N827, N819, N632, N756, N281);
nand NAND4 (N828, N826, N285, N140, N188);
and AND4 (N829, N809, N732, N399, N25);
xor XOR2 (N830, N807, N157);
nor NOR3 (N831, N823, N74, N374);
nor NOR2 (N832, N827, N469);
not NOT1 (N833, N830);
xor XOR2 (N834, N815, N822);
and AND4 (N835, N828, N609, N345, N805);
or OR2 (N836, N780, N150);
buf BUF1 (N837, N825);
buf BUF1 (N838, N837);
xor XOR2 (N839, N833, N634);
not NOT1 (N840, N836);
and AND3 (N841, N839, N275, N699);
nand NAND4 (N842, N840, N726, N217, N706);
buf BUF1 (N843, N832);
nor NOR2 (N844, N831, N218);
nor NOR4 (N845, N829, N783, N382, N579);
xor XOR2 (N846, N844, N756);
xor XOR2 (N847, N845, N154);
nand NAND3 (N848, N842, N275, N301);
xor XOR2 (N849, N846, N385);
nand NAND2 (N850, N838, N524);
not NOT1 (N851, N817);
buf BUF1 (N852, N849);
not NOT1 (N853, N835);
or OR4 (N854, N843, N639, N520, N295);
nand NAND2 (N855, N854, N552);
not NOT1 (N856, N852);
or OR2 (N857, N855, N850);
not NOT1 (N858, N356);
buf BUF1 (N859, N856);
xor XOR2 (N860, N858, N618);
nor NOR2 (N861, N853, N693);
nor NOR2 (N862, N848, N748);
and AND3 (N863, N857, N858, N128);
or OR3 (N864, N860, N676, N404);
not NOT1 (N865, N861);
buf BUF1 (N866, N865);
or OR3 (N867, N863, N511, N692);
xor XOR2 (N868, N862, N711);
nand NAND4 (N869, N868, N808, N44, N841);
buf BUF1 (N870, N158);
not NOT1 (N871, N847);
nor NOR3 (N872, N820, N483, N344);
nand NAND4 (N873, N869, N225, N522, N551);
nand NAND4 (N874, N870, N92, N27, N63);
xor XOR2 (N875, N866, N125);
or OR3 (N876, N864, N473, N407);
and AND2 (N877, N876, N809);
buf BUF1 (N878, N873);
and AND2 (N879, N878, N311);
xor XOR2 (N880, N867, N579);
and AND2 (N881, N875, N30);
buf BUF1 (N882, N871);
buf BUF1 (N883, N872);
nor NOR2 (N884, N879, N352);
and AND4 (N885, N884, N138, N164, N288);
not NOT1 (N886, N880);
xor XOR2 (N887, N886, N29);
xor XOR2 (N888, N883, N353);
xor XOR2 (N889, N885, N730);
buf BUF1 (N890, N851);
nand NAND2 (N891, N890, N699);
or OR4 (N892, N834, N301, N890, N158);
and AND3 (N893, N874, N82, N328);
buf BUF1 (N894, N859);
buf BUF1 (N895, N892);
nand NAND4 (N896, N882, N12, N429, N556);
nand NAND2 (N897, N891, N171);
not NOT1 (N898, N887);
nand NAND3 (N899, N881, N234, N216);
xor XOR2 (N900, N893, N849);
not NOT1 (N901, N898);
nand NAND3 (N902, N899, N716, N128);
and AND4 (N903, N902, N868, N160, N456);
or OR2 (N904, N903, N626);
not NOT1 (N905, N904);
and AND3 (N906, N889, N700, N705);
and AND2 (N907, N905, N342);
or OR4 (N908, N896, N98, N280, N299);
xor XOR2 (N909, N900, N242);
nand NAND3 (N910, N908, N569, N103);
and AND2 (N911, N910, N86);
buf BUF1 (N912, N911);
nand NAND2 (N913, N895, N96);
xor XOR2 (N914, N913, N171);
and AND3 (N915, N909, N68, N164);
nor NOR3 (N916, N901, N833, N896);
or OR2 (N917, N916, N570);
nor NOR3 (N918, N906, N585, N244);
or OR4 (N919, N894, N391, N538, N315);
nand NAND2 (N920, N915, N2);
or OR3 (N921, N917, N64, N743);
xor XOR2 (N922, N888, N873);
nand NAND2 (N923, N918, N525);
nand NAND3 (N924, N914, N459, N214);
nand NAND2 (N925, N922, N315);
nand NAND2 (N926, N919, N460);
or OR3 (N927, N912, N525, N577);
nor NOR3 (N928, N897, N121, N366);
buf BUF1 (N929, N907);
not NOT1 (N930, N928);
and AND4 (N931, N924, N745, N409, N785);
and AND4 (N932, N920, N917, N129, N635);
buf BUF1 (N933, N925);
nand NAND3 (N934, N921, N246, N902);
nand NAND2 (N935, N932, N345);
and AND3 (N936, N923, N393, N515);
nand NAND3 (N937, N926, N384, N218);
and AND3 (N938, N936, N127, N555);
not NOT1 (N939, N877);
and AND2 (N940, N937, N794);
xor XOR2 (N941, N934, N697);
nand NAND2 (N942, N930, N276);
xor XOR2 (N943, N940, N179);
nor NOR4 (N944, N942, N329, N352, N856);
nor NOR4 (N945, N939, N164, N865, N247);
or OR3 (N946, N929, N139, N492);
or OR2 (N947, N941, N27);
or OR3 (N948, N938, N858, N506);
buf BUF1 (N949, N935);
nor NOR4 (N950, N931, N279, N90, N601);
nor NOR4 (N951, N945, N493, N763, N760);
or OR3 (N952, N949, N130, N692);
nor NOR3 (N953, N946, N49, N609);
nor NOR3 (N954, N948, N550, N525);
nand NAND3 (N955, N947, N865, N99);
not NOT1 (N956, N943);
nand NAND2 (N957, N933, N278);
nor NOR4 (N958, N944, N484, N393, N529);
buf BUF1 (N959, N956);
nand NAND3 (N960, N952, N860, N126);
xor XOR2 (N961, N951, N123);
not NOT1 (N962, N957);
not NOT1 (N963, N958);
buf BUF1 (N964, N950);
buf BUF1 (N965, N963);
xor XOR2 (N966, N965, N792);
buf BUF1 (N967, N953);
nand NAND4 (N968, N954, N416, N602, N908);
nor NOR3 (N969, N967, N747, N325);
nor NOR2 (N970, N955, N903);
or OR3 (N971, N961, N160, N70);
buf BUF1 (N972, N966);
buf BUF1 (N973, N969);
nand NAND3 (N974, N964, N259, N334);
not NOT1 (N975, N960);
nand NAND4 (N976, N971, N268, N901, N362);
nor NOR2 (N977, N976, N944);
not NOT1 (N978, N973);
xor XOR2 (N979, N977, N74);
and AND2 (N980, N978, N394);
or OR4 (N981, N970, N498, N72, N603);
not NOT1 (N982, N968);
nor NOR2 (N983, N974, N190);
nand NAND4 (N984, N962, N401, N521, N180);
or OR4 (N985, N984, N958, N930, N677);
or OR2 (N986, N959, N678);
buf BUF1 (N987, N979);
nor NOR4 (N988, N975, N553, N164, N959);
nand NAND3 (N989, N985, N52, N113);
nand NAND3 (N990, N986, N956, N367);
nor NOR4 (N991, N983, N183, N130, N911);
nor NOR2 (N992, N990, N244);
xor XOR2 (N993, N980, N336);
and AND4 (N994, N972, N677, N556, N213);
nand NAND4 (N995, N981, N714, N236, N380);
not NOT1 (N996, N992);
xor XOR2 (N997, N988, N222);
and AND3 (N998, N927, N928, N565);
xor XOR2 (N999, N987, N950);
nand NAND3 (N1000, N996, N862, N269);
nor NOR3 (N1001, N982, N785, N768);
xor XOR2 (N1002, N1001, N799);
buf BUF1 (N1003, N994);
not NOT1 (N1004, N997);
xor XOR2 (N1005, N995, N543);
xor XOR2 (N1006, N1000, N30);
and AND4 (N1007, N998, N1004, N939, N608);
nor NOR2 (N1008, N430, N934);
nand NAND3 (N1009, N1002, N463, N649);
buf BUF1 (N1010, N993);
buf BUF1 (N1011, N1008);
xor XOR2 (N1012, N1006, N997);
nand NAND2 (N1013, N999, N814);
and AND4 (N1014, N1003, N645, N45, N281);
not NOT1 (N1015, N991);
xor XOR2 (N1016, N1015, N663);
not NOT1 (N1017, N1011);
nand NAND4 (N1018, N989, N347, N290, N768);
or OR4 (N1019, N1005, N543, N1, N377);
not NOT1 (N1020, N1019);
nor NOR3 (N1021, N1020, N1004, N263);
buf BUF1 (N1022, N1021);
nor NOR2 (N1023, N1017, N6);
nand NAND4 (N1024, N1012, N840, N163, N401);
nand NAND3 (N1025, N1023, N630, N242);
xor XOR2 (N1026, N1024, N715);
or OR4 (N1027, N1009, N7, N286, N158);
nand NAND2 (N1028, N1026, N118);
nand NAND4 (N1029, N1025, N293, N765, N651);
xor XOR2 (N1030, N1016, N452);
and AND2 (N1031, N1022, N434);
and AND2 (N1032, N1014, N740);
not NOT1 (N1033, N1031);
xor XOR2 (N1034, N1010, N532);
not NOT1 (N1035, N1018);
nor NOR4 (N1036, N1032, N717, N30, N705);
not NOT1 (N1037, N1027);
buf BUF1 (N1038, N1013);
nor NOR3 (N1039, N1028, N65, N618);
nor NOR2 (N1040, N1030, N238);
xor XOR2 (N1041, N1034, N326);
nor NOR2 (N1042, N1038, N493);
nand NAND3 (N1043, N1035, N483, N628);
xor XOR2 (N1044, N1041, N213);
xor XOR2 (N1045, N1029, N386);
nand NAND3 (N1046, N1044, N570, N52);
or OR3 (N1047, N1040, N613, N107);
buf BUF1 (N1048, N1033);
buf BUF1 (N1049, N1045);
and AND3 (N1050, N1039, N723, N17);
and AND3 (N1051, N1049, N960, N454);
and AND4 (N1052, N1007, N960, N255, N782);
or OR3 (N1053, N1042, N939, N885);
buf BUF1 (N1054, N1050);
buf BUF1 (N1055, N1051);
buf BUF1 (N1056, N1047);
nand NAND3 (N1057, N1053, N679, N585);
xor XOR2 (N1058, N1043, N977);
not NOT1 (N1059, N1048);
not NOT1 (N1060, N1055);
and AND4 (N1061, N1054, N451, N340, N475);
nor NOR3 (N1062, N1059, N30, N422);
buf BUF1 (N1063, N1060);
not NOT1 (N1064, N1036);
buf BUF1 (N1065, N1037);
or OR2 (N1066, N1063, N215);
not NOT1 (N1067, N1066);
buf BUF1 (N1068, N1058);
xor XOR2 (N1069, N1067, N1060);
and AND3 (N1070, N1065, N108, N695);
and AND4 (N1071, N1062, N420, N511, N838);
nor NOR2 (N1072, N1061, N60);
or OR2 (N1073, N1069, N146);
not NOT1 (N1074, N1052);
and AND4 (N1075, N1071, N189, N915, N1009);
and AND2 (N1076, N1073, N535);
buf BUF1 (N1077, N1070);
not NOT1 (N1078, N1056);
buf BUF1 (N1079, N1075);
or OR4 (N1080, N1072, N272, N424, N240);
and AND4 (N1081, N1074, N692, N367, N594);
xor XOR2 (N1082, N1046, N885);
nand NAND4 (N1083, N1077, N598, N496, N173);
not NOT1 (N1084, N1064);
nor NOR4 (N1085, N1076, N426, N537, N702);
nor NOR2 (N1086, N1079, N1075);
not NOT1 (N1087, N1068);
nand NAND2 (N1088, N1086, N734);
nand NAND2 (N1089, N1057, N662);
nor NOR2 (N1090, N1084, N862);
nor NOR4 (N1091, N1085, N121, N24, N633);
buf BUF1 (N1092, N1081);
or OR2 (N1093, N1088, N902);
and AND4 (N1094, N1082, N880, N303, N1032);
buf BUF1 (N1095, N1087);
buf BUF1 (N1096, N1089);
and AND2 (N1097, N1078, N101);
and AND4 (N1098, N1091, N749, N627, N299);
nor NOR2 (N1099, N1092, N469);
and AND2 (N1100, N1093, N478);
xor XOR2 (N1101, N1097, N472);
buf BUF1 (N1102, N1094);
and AND3 (N1103, N1080, N569, N104);
and AND4 (N1104, N1103, N836, N72, N347);
or OR2 (N1105, N1083, N205);
nand NAND3 (N1106, N1100, N270, N1096);
not NOT1 (N1107, N199);
nor NOR3 (N1108, N1090, N27, N765);
or OR3 (N1109, N1105, N553, N797);
nor NOR2 (N1110, N1106, N68);
xor XOR2 (N1111, N1098, N109);
xor XOR2 (N1112, N1110, N764);
xor XOR2 (N1113, N1102, N822);
buf BUF1 (N1114, N1109);
not NOT1 (N1115, N1108);
nor NOR2 (N1116, N1113, N1073);
or OR2 (N1117, N1095, N527);
nand NAND4 (N1118, N1111, N780, N441, N760);
xor XOR2 (N1119, N1114, N801);
nor NOR2 (N1120, N1099, N913);
nor NOR3 (N1121, N1115, N51, N179);
xor XOR2 (N1122, N1107, N334);
or OR3 (N1123, N1120, N742, N463);
buf BUF1 (N1124, N1121);
and AND3 (N1125, N1123, N752, N393);
buf BUF1 (N1126, N1101);
nand NAND3 (N1127, N1118, N658, N193);
buf BUF1 (N1128, N1124);
xor XOR2 (N1129, N1125, N352);
and AND4 (N1130, N1104, N817, N191, N1122);
xor XOR2 (N1131, N468, N781);
xor XOR2 (N1132, N1130, N279);
or OR4 (N1133, N1132, N1060, N440, N371);
nor NOR4 (N1134, N1129, N816, N984, N956);
xor XOR2 (N1135, N1117, N738);
xor XOR2 (N1136, N1127, N425);
nor NOR2 (N1137, N1134, N937);
buf BUF1 (N1138, N1131);
xor XOR2 (N1139, N1135, N489);
not NOT1 (N1140, N1126);
xor XOR2 (N1141, N1133, N103);
and AND2 (N1142, N1138, N26);
and AND3 (N1143, N1116, N328, N56);
nor NOR3 (N1144, N1112, N311, N9);
and AND3 (N1145, N1140, N932, N757);
and AND4 (N1146, N1136, N216, N1037, N757);
nor NOR3 (N1147, N1141, N139, N141);
nand NAND2 (N1148, N1137, N133);
or OR4 (N1149, N1128, N993, N498, N58);
not NOT1 (N1150, N1142);
buf BUF1 (N1151, N1145);
and AND3 (N1152, N1144, N738, N102);
buf BUF1 (N1153, N1152);
buf BUF1 (N1154, N1153);
or OR3 (N1155, N1148, N885, N471);
nor NOR4 (N1156, N1149, N853, N121, N49);
nor NOR3 (N1157, N1147, N1136, N890);
nor NOR3 (N1158, N1155, N82, N305);
buf BUF1 (N1159, N1119);
nor NOR2 (N1160, N1156, N1089);
buf BUF1 (N1161, N1139);
or OR2 (N1162, N1143, N1072);
and AND4 (N1163, N1159, N550, N545, N942);
buf BUF1 (N1164, N1162);
xor XOR2 (N1165, N1146, N248);
nor NOR3 (N1166, N1161, N562, N1052);
buf BUF1 (N1167, N1157);
buf BUF1 (N1168, N1158);
not NOT1 (N1169, N1150);
and AND4 (N1170, N1163, N1074, N1026, N312);
and AND2 (N1171, N1169, N1073);
not NOT1 (N1172, N1165);
xor XOR2 (N1173, N1160, N37);
not NOT1 (N1174, N1171);
or OR3 (N1175, N1168, N1134, N1050);
not NOT1 (N1176, N1164);
and AND3 (N1177, N1170, N730, N289);
buf BUF1 (N1178, N1166);
xor XOR2 (N1179, N1177, N1162);
xor XOR2 (N1180, N1154, N1046);
not NOT1 (N1181, N1175);
nand NAND2 (N1182, N1176, N650);
nor NOR3 (N1183, N1181, N553, N1178);
xor XOR2 (N1184, N762, N638);
buf BUF1 (N1185, N1184);
not NOT1 (N1186, N1151);
and AND3 (N1187, N1173, N54, N95);
nor NOR4 (N1188, N1185, N229, N305, N7);
not NOT1 (N1189, N1172);
and AND4 (N1190, N1183, N311, N576, N857);
nand NAND2 (N1191, N1179, N508);
nor NOR3 (N1192, N1190, N571, N1050);
nand NAND2 (N1193, N1174, N1002);
nand NAND2 (N1194, N1192, N355);
not NOT1 (N1195, N1186);
not NOT1 (N1196, N1182);
not NOT1 (N1197, N1187);
or OR2 (N1198, N1167, N673);
nor NOR4 (N1199, N1195, N1050, N995, N599);
xor XOR2 (N1200, N1191, N222);
xor XOR2 (N1201, N1189, N513);
not NOT1 (N1202, N1196);
xor XOR2 (N1203, N1180, N575);
buf BUF1 (N1204, N1199);
not NOT1 (N1205, N1201);
and AND4 (N1206, N1193, N1199, N1157, N34);
nor NOR4 (N1207, N1204, N578, N642, N123);
nand NAND2 (N1208, N1194, N33);
nor NOR4 (N1209, N1200, N838, N109, N595);
buf BUF1 (N1210, N1205);
nand NAND4 (N1211, N1207, N467, N1000, N22);
or OR3 (N1212, N1198, N657, N731);
nand NAND3 (N1213, N1203, N196, N241);
or OR2 (N1214, N1197, N814);
nor NOR4 (N1215, N1202, N403, N1158, N606);
nor NOR3 (N1216, N1212, N924, N762);
not NOT1 (N1217, N1215);
nor NOR4 (N1218, N1214, N88, N696, N822);
nand NAND4 (N1219, N1188, N568, N622, N1016);
or OR3 (N1220, N1216, N626, N858);
buf BUF1 (N1221, N1220);
not NOT1 (N1222, N1211);
not NOT1 (N1223, N1213);
xor XOR2 (N1224, N1219, N277);
and AND4 (N1225, N1206, N674, N98, N1116);
buf BUF1 (N1226, N1218);
xor XOR2 (N1227, N1221, N78);
not NOT1 (N1228, N1227);
not NOT1 (N1229, N1222);
and AND4 (N1230, N1224, N209, N349, N456);
nor NOR2 (N1231, N1229, N1030);
and AND2 (N1232, N1228, N46);
nand NAND4 (N1233, N1225, N195, N66, N31);
and AND4 (N1234, N1233, N418, N801, N663);
nand NAND3 (N1235, N1223, N337, N188);
nand NAND4 (N1236, N1232, N1157, N703, N966);
buf BUF1 (N1237, N1217);
nand NAND2 (N1238, N1210, N588);
nand NAND4 (N1239, N1238, N884, N863, N375);
buf BUF1 (N1240, N1226);
or OR2 (N1241, N1235, N148);
xor XOR2 (N1242, N1236, N584);
buf BUF1 (N1243, N1237);
nor NOR2 (N1244, N1243, N326);
not NOT1 (N1245, N1209);
or OR3 (N1246, N1234, N898, N328);
nor NOR2 (N1247, N1231, N808);
or OR2 (N1248, N1208, N878);
or OR2 (N1249, N1246, N159);
nor NOR2 (N1250, N1244, N1060);
and AND2 (N1251, N1242, N910);
not NOT1 (N1252, N1250);
or OR2 (N1253, N1251, N26);
xor XOR2 (N1254, N1253, N74);
and AND2 (N1255, N1249, N9);
xor XOR2 (N1256, N1247, N247);
and AND2 (N1257, N1240, N1028);
nand NAND2 (N1258, N1239, N92);
buf BUF1 (N1259, N1258);
or OR2 (N1260, N1241, N873);
nor NOR2 (N1261, N1248, N922);
nor NOR2 (N1262, N1245, N106);
nand NAND3 (N1263, N1252, N467, N606);
or OR3 (N1264, N1260, N978, N245);
and AND2 (N1265, N1256, N728);
and AND4 (N1266, N1259, N418, N659, N818);
nand NAND3 (N1267, N1255, N302, N65);
nor NOR2 (N1268, N1230, N736);
and AND4 (N1269, N1263, N642, N673, N165);
or OR4 (N1270, N1264, N1135, N109, N1127);
and AND2 (N1271, N1257, N852);
or OR4 (N1272, N1254, N1113, N1089, N330);
xor XOR2 (N1273, N1266, N1217);
xor XOR2 (N1274, N1267, N252);
or OR3 (N1275, N1269, N852, N625);
xor XOR2 (N1276, N1261, N795);
nand NAND2 (N1277, N1268, N538);
buf BUF1 (N1278, N1275);
buf BUF1 (N1279, N1277);
nand NAND2 (N1280, N1271, N738);
xor XOR2 (N1281, N1280, N865);
buf BUF1 (N1282, N1281);
buf BUF1 (N1283, N1278);
nand NAND4 (N1284, N1276, N59, N887, N1226);
and AND2 (N1285, N1283, N992);
and AND4 (N1286, N1274, N219, N439, N265);
or OR4 (N1287, N1265, N976, N568, N776);
and AND2 (N1288, N1270, N23);
and AND3 (N1289, N1287, N257, N348);
buf BUF1 (N1290, N1282);
buf BUF1 (N1291, N1286);
buf BUF1 (N1292, N1290);
nand NAND2 (N1293, N1291, N605);
xor XOR2 (N1294, N1288, N921);
xor XOR2 (N1295, N1292, N1180);
buf BUF1 (N1296, N1284);
xor XOR2 (N1297, N1262, N93);
or OR3 (N1298, N1272, N984, N550);
or OR2 (N1299, N1296, N512);
nand NAND4 (N1300, N1297, N79, N72, N815);
not NOT1 (N1301, N1289);
nand NAND2 (N1302, N1285, N235);
buf BUF1 (N1303, N1301);
buf BUF1 (N1304, N1302);
or OR3 (N1305, N1279, N902, N699);
or OR4 (N1306, N1299, N1219, N975, N1156);
or OR3 (N1307, N1298, N983, N395);
buf BUF1 (N1308, N1273);
xor XOR2 (N1309, N1294, N14);
or OR3 (N1310, N1304, N1246, N178);
not NOT1 (N1311, N1310);
nand NAND3 (N1312, N1293, N1102, N733);
nand NAND2 (N1313, N1312, N113);
nand NAND4 (N1314, N1306, N23, N348, N384);
or OR3 (N1315, N1305, N101, N1025);
or OR2 (N1316, N1311, N953);
or OR2 (N1317, N1300, N284);
and AND2 (N1318, N1316, N312);
buf BUF1 (N1319, N1308);
buf BUF1 (N1320, N1309);
nand NAND2 (N1321, N1315, N656);
and AND3 (N1322, N1317, N1304, N417);
or OR3 (N1323, N1313, N567, N213);
xor XOR2 (N1324, N1295, N1141);
not NOT1 (N1325, N1320);
nor NOR2 (N1326, N1307, N941);
buf BUF1 (N1327, N1323);
buf BUF1 (N1328, N1325);
and AND3 (N1329, N1303, N850, N1054);
nand NAND2 (N1330, N1322, N888);
and AND2 (N1331, N1330, N236);
buf BUF1 (N1332, N1329);
buf BUF1 (N1333, N1319);
and AND3 (N1334, N1326, N211, N108);
xor XOR2 (N1335, N1318, N313);
xor XOR2 (N1336, N1324, N1165);
xor XOR2 (N1337, N1336, N1037);
not NOT1 (N1338, N1314);
buf BUF1 (N1339, N1327);
xor XOR2 (N1340, N1337, N309);
or OR4 (N1341, N1340, N1241, N136, N1256);
nor NOR3 (N1342, N1332, N749, N74);
nor NOR4 (N1343, N1338, N536, N306, N749);
and AND4 (N1344, N1342, N1268, N763, N1116);
xor XOR2 (N1345, N1321, N69);
and AND2 (N1346, N1345, N328);
and AND3 (N1347, N1341, N608, N649);
not NOT1 (N1348, N1331);
xor XOR2 (N1349, N1334, N445);
and AND3 (N1350, N1343, N49, N211);
and AND4 (N1351, N1335, N97, N1305, N731);
xor XOR2 (N1352, N1346, N1089);
xor XOR2 (N1353, N1352, N1080);
buf BUF1 (N1354, N1347);
not NOT1 (N1355, N1353);
buf BUF1 (N1356, N1348);
or OR3 (N1357, N1356, N2, N143);
nor NOR4 (N1358, N1333, N709, N927, N862);
nor NOR3 (N1359, N1328, N628, N199);
nor NOR4 (N1360, N1354, N1264, N1259, N382);
not NOT1 (N1361, N1350);
buf BUF1 (N1362, N1358);
not NOT1 (N1363, N1349);
not NOT1 (N1364, N1363);
or OR3 (N1365, N1355, N863, N730);
and AND4 (N1366, N1361, N960, N775, N1210);
nand NAND4 (N1367, N1360, N188, N1007, N1061);
nand NAND2 (N1368, N1362, N140);
nor NOR4 (N1369, N1365, N356, N660, N317);
buf BUF1 (N1370, N1369);
nor NOR2 (N1371, N1364, N191);
nor NOR2 (N1372, N1368, N820);
or OR2 (N1373, N1344, N360);
not NOT1 (N1374, N1351);
nor NOR4 (N1375, N1359, N1019, N826, N824);
buf BUF1 (N1376, N1372);
or OR3 (N1377, N1366, N781, N763);
buf BUF1 (N1378, N1373);
buf BUF1 (N1379, N1378);
or OR2 (N1380, N1379, N554);
xor XOR2 (N1381, N1339, N617);
and AND2 (N1382, N1381, N375);
not NOT1 (N1383, N1375);
and AND3 (N1384, N1370, N1102, N690);
not NOT1 (N1385, N1357);
buf BUF1 (N1386, N1383);
xor XOR2 (N1387, N1377, N1086);
nor NOR2 (N1388, N1387, N1156);
or OR3 (N1389, N1374, N1256, N385);
buf BUF1 (N1390, N1380);
and AND3 (N1391, N1386, N645, N483);
nand NAND3 (N1392, N1382, N102, N920);
nor NOR4 (N1393, N1389, N831, N797, N1064);
not NOT1 (N1394, N1367);
or OR3 (N1395, N1391, N6, N1062);
buf BUF1 (N1396, N1394);
nor NOR4 (N1397, N1392, N50, N1287, N131);
or OR3 (N1398, N1397, N1354, N1166);
xor XOR2 (N1399, N1385, N214);
nor NOR4 (N1400, N1390, N268, N243, N1088);
xor XOR2 (N1401, N1398, N311);
nand NAND4 (N1402, N1376, N145, N1257, N920);
nor NOR2 (N1403, N1396, N148);
nor NOR3 (N1404, N1400, N87, N105);
nand NAND3 (N1405, N1404, N784, N545);
nor NOR2 (N1406, N1384, N506);
nor NOR3 (N1407, N1395, N987, N185);
and AND3 (N1408, N1371, N1177, N774);
or OR4 (N1409, N1406, N1330, N1179, N1196);
nand NAND4 (N1410, N1388, N553, N430, N282);
xor XOR2 (N1411, N1399, N12);
and AND2 (N1412, N1401, N156);
nor NOR3 (N1413, N1412, N965, N201);
not NOT1 (N1414, N1410);
nand NAND2 (N1415, N1413, N646);
and AND4 (N1416, N1405, N686, N616, N86);
nor NOR4 (N1417, N1414, N410, N908, N3);
nor NOR4 (N1418, N1393, N1142, N782, N736);
nand NAND3 (N1419, N1415, N330, N856);
and AND4 (N1420, N1419, N428, N515, N748);
or OR3 (N1421, N1417, N1050, N1162);
or OR4 (N1422, N1402, N300, N1263, N133);
buf BUF1 (N1423, N1420);
xor XOR2 (N1424, N1407, N712);
xor XOR2 (N1425, N1421, N149);
xor XOR2 (N1426, N1423, N1059);
xor XOR2 (N1427, N1408, N1397);
and AND2 (N1428, N1422, N348);
xor XOR2 (N1429, N1424, N150);
buf BUF1 (N1430, N1428);
and AND2 (N1431, N1411, N605);
not NOT1 (N1432, N1416);
nand NAND3 (N1433, N1403, N1344, N532);
xor XOR2 (N1434, N1409, N539);
nand NAND2 (N1435, N1430, N213);
nand NAND4 (N1436, N1425, N34, N849, N97);
and AND2 (N1437, N1426, N52);
xor XOR2 (N1438, N1429, N580);
nand NAND4 (N1439, N1433, N1296, N152, N452);
not NOT1 (N1440, N1438);
and AND2 (N1441, N1436, N1186);
and AND3 (N1442, N1440, N1392, N348);
nand NAND4 (N1443, N1434, N1417, N1004, N342);
nand NAND4 (N1444, N1431, N650, N468, N396);
not NOT1 (N1445, N1443);
or OR3 (N1446, N1439, N1197, N1388);
and AND4 (N1447, N1444, N1120, N1063, N518);
xor XOR2 (N1448, N1441, N516);
nor NOR3 (N1449, N1448, N26, N1063);
buf BUF1 (N1450, N1449);
buf BUF1 (N1451, N1442);
buf BUF1 (N1452, N1437);
buf BUF1 (N1453, N1432);
and AND2 (N1454, N1427, N66);
nor NOR4 (N1455, N1447, N256, N460, N720);
or OR4 (N1456, N1435, N121, N172, N185);
not NOT1 (N1457, N1450);
buf BUF1 (N1458, N1445);
nand NAND2 (N1459, N1451, N758);
nor NOR3 (N1460, N1456, N221, N201);
xor XOR2 (N1461, N1460, N861);
and AND2 (N1462, N1454, N495);
nand NAND2 (N1463, N1459, N1144);
buf BUF1 (N1464, N1458);
xor XOR2 (N1465, N1463, N406);
buf BUF1 (N1466, N1465);
not NOT1 (N1467, N1462);
xor XOR2 (N1468, N1467, N168);
or OR2 (N1469, N1452, N351);
buf BUF1 (N1470, N1468);
or OR2 (N1471, N1453, N455);
nand NAND3 (N1472, N1457, N1091, N577);
nand NAND4 (N1473, N1470, N1344, N729, N968);
xor XOR2 (N1474, N1471, N972);
buf BUF1 (N1475, N1472);
and AND3 (N1476, N1466, N662, N609);
not NOT1 (N1477, N1475);
xor XOR2 (N1478, N1418, N404);
nand NAND3 (N1479, N1473, N639, N1110);
nand NAND3 (N1480, N1469, N1401, N1347);
and AND4 (N1481, N1477, N1315, N974, N248);
buf BUF1 (N1482, N1479);
or OR4 (N1483, N1482, N481, N75, N903);
buf BUF1 (N1484, N1461);
or OR2 (N1485, N1481, N717);
not NOT1 (N1486, N1474);
xor XOR2 (N1487, N1464, N886);
nor NOR4 (N1488, N1480, N514, N1240, N957);
or OR2 (N1489, N1455, N1168);
nor NOR2 (N1490, N1485, N587);
xor XOR2 (N1491, N1486, N449);
buf BUF1 (N1492, N1446);
not NOT1 (N1493, N1492);
nand NAND3 (N1494, N1490, N439, N996);
buf BUF1 (N1495, N1476);
buf BUF1 (N1496, N1491);
xor XOR2 (N1497, N1478, N1382);
nor NOR4 (N1498, N1489, N636, N551, N820);
or OR3 (N1499, N1487, N134, N1041);
xor XOR2 (N1500, N1488, N593);
xor XOR2 (N1501, N1483, N1182);
xor XOR2 (N1502, N1499, N785);
or OR3 (N1503, N1495, N1234, N418);
not NOT1 (N1504, N1500);
nand NAND3 (N1505, N1498, N1215, N148);
nand NAND3 (N1506, N1501, N764, N1344);
not NOT1 (N1507, N1506);
not NOT1 (N1508, N1493);
not NOT1 (N1509, N1496);
buf BUF1 (N1510, N1494);
or OR2 (N1511, N1503, N1246);
xor XOR2 (N1512, N1504, N636);
and AND4 (N1513, N1510, N725, N1350, N442);
or OR3 (N1514, N1509, N144, N657);
nand NAND4 (N1515, N1507, N1152, N82, N715);
xor XOR2 (N1516, N1513, N951);
or OR4 (N1517, N1502, N964, N127, N1190);
or OR2 (N1518, N1511, N731);
xor XOR2 (N1519, N1518, N32);
or OR2 (N1520, N1484, N622);
buf BUF1 (N1521, N1508);
nor NOR2 (N1522, N1515, N875);
xor XOR2 (N1523, N1521, N741);
nor NOR4 (N1524, N1522, N2, N559, N497);
nor NOR3 (N1525, N1512, N212, N28);
nand NAND3 (N1526, N1523, N601, N856);
xor XOR2 (N1527, N1526, N847);
buf BUF1 (N1528, N1514);
nand NAND3 (N1529, N1525, N428, N213);
nand NAND2 (N1530, N1520, N52);
buf BUF1 (N1531, N1529);
or OR4 (N1532, N1497, N934, N1361, N1289);
and AND2 (N1533, N1531, N660);
buf BUF1 (N1534, N1533);
and AND3 (N1535, N1519, N1301, N893);
nor NOR3 (N1536, N1532, N1155, N1202);
not NOT1 (N1537, N1527);
and AND4 (N1538, N1536, N386, N128, N1208);
or OR4 (N1539, N1537, N670, N260, N969);
not NOT1 (N1540, N1505);
xor XOR2 (N1541, N1530, N406);
buf BUF1 (N1542, N1540);
nand NAND4 (N1543, N1542, N123, N1064, N361);
and AND4 (N1544, N1538, N549, N196, N620);
nor NOR3 (N1545, N1541, N595, N528);
or OR3 (N1546, N1534, N720, N736);
buf BUF1 (N1547, N1544);
xor XOR2 (N1548, N1524, N1093);
nand NAND2 (N1549, N1539, N639);
not NOT1 (N1550, N1547);
nor NOR4 (N1551, N1535, N361, N215, N1041);
or OR4 (N1552, N1543, N797, N439, N1425);
and AND4 (N1553, N1545, N1535, N1477, N1102);
nand NAND2 (N1554, N1516, N734);
nor NOR2 (N1555, N1550, N1267);
or OR2 (N1556, N1548, N783);
buf BUF1 (N1557, N1556);
nor NOR3 (N1558, N1553, N673, N621);
and AND3 (N1559, N1552, N1354, N216);
buf BUF1 (N1560, N1517);
not NOT1 (N1561, N1560);
not NOT1 (N1562, N1559);
or OR3 (N1563, N1561, N1219, N1351);
buf BUF1 (N1564, N1528);
nor NOR3 (N1565, N1564, N756, N13);
buf BUF1 (N1566, N1563);
and AND4 (N1567, N1554, N1275, N784, N628);
nor NOR4 (N1568, N1558, N616, N738, N721);
or OR2 (N1569, N1551, N109);
buf BUF1 (N1570, N1555);
nor NOR3 (N1571, N1568, N1367, N492);
nor NOR4 (N1572, N1567, N388, N518, N1035);
and AND3 (N1573, N1572, N1191, N1069);
xor XOR2 (N1574, N1549, N121);
and AND4 (N1575, N1557, N73, N932, N1367);
nor NOR3 (N1576, N1546, N567, N428);
not NOT1 (N1577, N1565);
and AND3 (N1578, N1574, N1377, N471);
buf BUF1 (N1579, N1573);
and AND2 (N1580, N1575, N172);
xor XOR2 (N1581, N1570, N419);
xor XOR2 (N1582, N1580, N77);
buf BUF1 (N1583, N1571);
nor NOR4 (N1584, N1566, N41, N74, N503);
xor XOR2 (N1585, N1577, N158);
nand NAND4 (N1586, N1576, N1113, N299, N461);
and AND4 (N1587, N1578, N426, N177, N1099);
not NOT1 (N1588, N1584);
not NOT1 (N1589, N1581);
not NOT1 (N1590, N1586);
buf BUF1 (N1591, N1589);
nor NOR3 (N1592, N1588, N1168, N360);
buf BUF1 (N1593, N1591);
nand NAND2 (N1594, N1582, N1013);
nand NAND3 (N1595, N1562, N1443, N533);
buf BUF1 (N1596, N1585);
buf BUF1 (N1597, N1587);
buf BUF1 (N1598, N1590);
nor NOR3 (N1599, N1569, N1074, N1204);
or OR4 (N1600, N1594, N1275, N815, N74);
or OR3 (N1601, N1579, N1499, N817);
and AND4 (N1602, N1595, N295, N184, N818);
or OR2 (N1603, N1601, N371);
not NOT1 (N1604, N1592);
xor XOR2 (N1605, N1583, N1386);
and AND4 (N1606, N1597, N997, N470, N1532);
buf BUF1 (N1607, N1598);
buf BUF1 (N1608, N1603);
xor XOR2 (N1609, N1606, N1265);
nand NAND3 (N1610, N1593, N612, N1375);
nor NOR2 (N1611, N1608, N54);
and AND4 (N1612, N1605, N1101, N1454, N728);
xor XOR2 (N1613, N1596, N1080);
nor NOR4 (N1614, N1602, N577, N1014, N131);
and AND4 (N1615, N1610, N30, N1470, N367);
nor NOR3 (N1616, N1613, N549, N268);
nand NAND4 (N1617, N1615, N133, N1508, N690);
nor NOR2 (N1618, N1600, N419);
buf BUF1 (N1619, N1612);
nand NAND4 (N1620, N1616, N112, N39, N355);
nand NAND3 (N1621, N1618, N594, N1578);
or OR4 (N1622, N1604, N263, N518, N414);
or OR2 (N1623, N1609, N714);
nand NAND4 (N1624, N1614, N939, N1329, N1508);
nor NOR2 (N1625, N1621, N587);
xor XOR2 (N1626, N1623, N363);
and AND3 (N1627, N1622, N1163, N1011);
not NOT1 (N1628, N1626);
nand NAND3 (N1629, N1619, N1063, N450);
not NOT1 (N1630, N1607);
nor NOR4 (N1631, N1630, N459, N1077, N1472);
xor XOR2 (N1632, N1620, N650);
or OR4 (N1633, N1625, N1000, N1500, N825);
not NOT1 (N1634, N1628);
xor XOR2 (N1635, N1633, N46);
xor XOR2 (N1636, N1599, N1399);
nor NOR3 (N1637, N1611, N1448, N938);
nand NAND2 (N1638, N1635, N308);
buf BUF1 (N1639, N1638);
nor NOR2 (N1640, N1631, N698);
nand NAND2 (N1641, N1629, N754);
and AND3 (N1642, N1627, N330, N380);
nand NAND2 (N1643, N1617, N333);
buf BUF1 (N1644, N1639);
or OR3 (N1645, N1642, N1045, N1352);
xor XOR2 (N1646, N1644, N840);
buf BUF1 (N1647, N1646);
xor XOR2 (N1648, N1641, N1240);
nor NOR2 (N1649, N1636, N381);
xor XOR2 (N1650, N1647, N1062);
nand NAND3 (N1651, N1649, N568, N1337);
not NOT1 (N1652, N1650);
nor NOR3 (N1653, N1632, N1017, N1361);
xor XOR2 (N1654, N1653, N922);
xor XOR2 (N1655, N1643, N109);
or OR3 (N1656, N1634, N1113, N994);
buf BUF1 (N1657, N1656);
or OR2 (N1658, N1645, N1429);
and AND2 (N1659, N1624, N629);
not NOT1 (N1660, N1655);
and AND4 (N1661, N1659, N1365, N613, N189);
nand NAND3 (N1662, N1637, N1421, N213);
nor NOR3 (N1663, N1648, N1652, N1032);
or OR2 (N1664, N834, N483);
nand NAND3 (N1665, N1664, N881, N1503);
xor XOR2 (N1666, N1662, N461);
nand NAND4 (N1667, N1665, N1493, N1413, N769);
xor XOR2 (N1668, N1654, N488);
or OR3 (N1669, N1660, N1385, N1505);
and AND2 (N1670, N1661, N1060);
nor NOR3 (N1671, N1667, N184, N1458);
nand NAND4 (N1672, N1651, N1059, N1183, N1070);
nor NOR4 (N1673, N1663, N420, N382, N244);
nor NOR2 (N1674, N1672, N1653);
nor NOR3 (N1675, N1669, N1420, N1391);
buf BUF1 (N1676, N1668);
xor XOR2 (N1677, N1666, N934);
buf BUF1 (N1678, N1673);
or OR3 (N1679, N1671, N1140, N208);
or OR3 (N1680, N1677, N979, N1572);
and AND2 (N1681, N1679, N555);
buf BUF1 (N1682, N1640);
buf BUF1 (N1683, N1676);
and AND2 (N1684, N1657, N928);
or OR2 (N1685, N1684, N1612);
not NOT1 (N1686, N1658);
or OR3 (N1687, N1674, N546, N1534);
not NOT1 (N1688, N1670);
buf BUF1 (N1689, N1686);
nor NOR3 (N1690, N1683, N69, N772);
nor NOR4 (N1691, N1675, N521, N1611, N546);
not NOT1 (N1692, N1685);
nor NOR3 (N1693, N1681, N44, N1659);
nand NAND4 (N1694, N1678, N1585, N203, N1302);
xor XOR2 (N1695, N1680, N458);
xor XOR2 (N1696, N1694, N1487);
buf BUF1 (N1697, N1692);
or OR2 (N1698, N1697, N428);
nor NOR4 (N1699, N1682, N1097, N1679, N811);
nor NOR3 (N1700, N1699, N1211, N848);
nand NAND4 (N1701, N1698, N810, N1459, N930);
not NOT1 (N1702, N1700);
nor NOR3 (N1703, N1693, N1103, N543);
buf BUF1 (N1704, N1689);
not NOT1 (N1705, N1703);
or OR3 (N1706, N1705, N283, N574);
buf BUF1 (N1707, N1688);
nor NOR2 (N1708, N1702, N986);
or OR4 (N1709, N1701, N561, N1200, N884);
xor XOR2 (N1710, N1690, N896);
nor NOR2 (N1711, N1691, N739);
or OR4 (N1712, N1711, N251, N676, N1308);
not NOT1 (N1713, N1712);
nand NAND3 (N1714, N1713, N819, N912);
and AND4 (N1715, N1687, N1327, N1399, N1312);
buf BUF1 (N1716, N1709);
nor NOR2 (N1717, N1695, N1074);
nand NAND2 (N1718, N1717, N373);
nand NAND3 (N1719, N1696, N1452, N161);
nand NAND4 (N1720, N1707, N104, N18, N478);
not NOT1 (N1721, N1719);
nand NAND2 (N1722, N1720, N1);
nand NAND2 (N1723, N1710, N394);
nand NAND3 (N1724, N1714, N1633, N245);
nor NOR4 (N1725, N1716, N1378, N1075, N1226);
nor NOR3 (N1726, N1723, N1619, N512);
or OR2 (N1727, N1706, N366);
not NOT1 (N1728, N1715);
xor XOR2 (N1729, N1721, N1726);
xor XOR2 (N1730, N1101, N385);
and AND4 (N1731, N1722, N1504, N969, N638);
not NOT1 (N1732, N1718);
nor NOR2 (N1733, N1708, N215);
nand NAND2 (N1734, N1733, N1490);
not NOT1 (N1735, N1727);
buf BUF1 (N1736, N1728);
xor XOR2 (N1737, N1732, N68);
buf BUF1 (N1738, N1736);
not NOT1 (N1739, N1729);
xor XOR2 (N1740, N1724, N17);
or OR4 (N1741, N1734, N1642, N1496, N943);
nand NAND2 (N1742, N1737, N1229);
or OR2 (N1743, N1741, N468);
xor XOR2 (N1744, N1725, N308);
and AND2 (N1745, N1738, N1296);
not NOT1 (N1746, N1743);
buf BUF1 (N1747, N1730);
nor NOR2 (N1748, N1704, N409);
nand NAND2 (N1749, N1748, N1152);
buf BUF1 (N1750, N1731);
and AND2 (N1751, N1744, N947);
nor NOR4 (N1752, N1739, N1256, N277, N12);
xor XOR2 (N1753, N1740, N1047);
nand NAND2 (N1754, N1735, N30);
xor XOR2 (N1755, N1746, N1468);
or OR3 (N1756, N1752, N416, N1392);
nor NOR2 (N1757, N1742, N1128);
xor XOR2 (N1758, N1757, N141);
nand NAND2 (N1759, N1753, N1014);
xor XOR2 (N1760, N1749, N513);
nor NOR2 (N1761, N1756, N891);
buf BUF1 (N1762, N1751);
not NOT1 (N1763, N1750);
and AND3 (N1764, N1754, N1420, N297);
nand NAND3 (N1765, N1760, N490, N37);
nor NOR2 (N1766, N1747, N427);
or OR4 (N1767, N1745, N718, N16, N1628);
not NOT1 (N1768, N1755);
nand NAND4 (N1769, N1764, N705, N1114, N928);
or OR3 (N1770, N1767, N760, N1114);
and AND2 (N1771, N1758, N1234);
not NOT1 (N1772, N1768);
not NOT1 (N1773, N1769);
not NOT1 (N1774, N1766);
nand NAND4 (N1775, N1772, N48, N162, N229);
nand NAND3 (N1776, N1765, N571, N975);
nand NAND2 (N1777, N1761, N1213);
nand NAND2 (N1778, N1774, N573);
nand NAND2 (N1779, N1771, N819);
xor XOR2 (N1780, N1778, N546);
nor NOR3 (N1781, N1780, N749, N1193);
not NOT1 (N1782, N1775);
nand NAND4 (N1783, N1781, N1778, N186, N155);
buf BUF1 (N1784, N1777);
nand NAND4 (N1785, N1770, N383, N540, N623);
and AND4 (N1786, N1763, N1661, N1276, N940);
nor NOR3 (N1787, N1762, N205, N1074);
and AND2 (N1788, N1784, N979);
and AND3 (N1789, N1759, N1202, N826);
and AND3 (N1790, N1776, N1756, N667);
xor XOR2 (N1791, N1787, N1723);
nor NOR3 (N1792, N1779, N59, N1658);
buf BUF1 (N1793, N1773);
and AND2 (N1794, N1786, N1142);
nor NOR2 (N1795, N1792, N460);
buf BUF1 (N1796, N1789);
or OR4 (N1797, N1796, N917, N1736, N1038);
xor XOR2 (N1798, N1797, N1451);
nor NOR2 (N1799, N1793, N784);
xor XOR2 (N1800, N1783, N650);
not NOT1 (N1801, N1791);
and AND3 (N1802, N1782, N1684, N77);
nor NOR3 (N1803, N1799, N654, N792);
and AND4 (N1804, N1795, N435, N67, N456);
xor XOR2 (N1805, N1794, N1089);
nor NOR4 (N1806, N1805, N1248, N956, N729);
or OR3 (N1807, N1802, N317, N327);
nor NOR3 (N1808, N1785, N211, N1413);
and AND3 (N1809, N1790, N810, N1287);
not NOT1 (N1810, N1798);
nor NOR3 (N1811, N1801, N745, N1034);
not NOT1 (N1812, N1807);
or OR3 (N1813, N1812, N784, N1478);
nand NAND3 (N1814, N1810, N724, N1540);
not NOT1 (N1815, N1804);
xor XOR2 (N1816, N1814, N1555);
nand NAND4 (N1817, N1803, N985, N690, N391);
or OR3 (N1818, N1788, N1529, N1443);
nor NOR3 (N1819, N1811, N1162, N455);
not NOT1 (N1820, N1819);
not NOT1 (N1821, N1813);
and AND3 (N1822, N1818, N1790, N434);
buf BUF1 (N1823, N1809);
buf BUF1 (N1824, N1817);
or OR3 (N1825, N1824, N1431, N720);
not NOT1 (N1826, N1823);
nand NAND2 (N1827, N1815, N1517);
buf BUF1 (N1828, N1821);
nand NAND4 (N1829, N1806, N1501, N48, N534);
nand NAND4 (N1830, N1816, N437, N833, N1382);
and AND2 (N1831, N1830, N858);
buf BUF1 (N1832, N1820);
nand NAND2 (N1833, N1825, N1521);
or OR2 (N1834, N1808, N1470);
buf BUF1 (N1835, N1827);
and AND2 (N1836, N1835, N1697);
xor XOR2 (N1837, N1831, N1692);
nor NOR3 (N1838, N1829, N832, N1239);
xor XOR2 (N1839, N1836, N1785);
xor XOR2 (N1840, N1800, N1250);
or OR4 (N1841, N1826, N291, N1366, N1453);
nand NAND3 (N1842, N1833, N1767, N110);
buf BUF1 (N1843, N1834);
nor NOR2 (N1844, N1828, N1373);
buf BUF1 (N1845, N1840);
and AND3 (N1846, N1838, N72, N66);
nand NAND4 (N1847, N1844, N697, N24, N157);
buf BUF1 (N1848, N1832);
nand NAND2 (N1849, N1837, N666);
xor XOR2 (N1850, N1847, N602);
or OR4 (N1851, N1845, N1180, N1333, N814);
nor NOR3 (N1852, N1851, N1776, N1509);
nor NOR3 (N1853, N1843, N1218, N1291);
and AND4 (N1854, N1842, N545, N159, N1254);
or OR2 (N1855, N1852, N408);
nor NOR3 (N1856, N1848, N620, N1424);
and AND2 (N1857, N1849, N566);
xor XOR2 (N1858, N1822, N513);
nor NOR4 (N1859, N1841, N55, N820, N157);
nor NOR4 (N1860, N1846, N968, N609, N507);
nand NAND4 (N1861, N1858, N502, N811, N1152);
or OR4 (N1862, N1850, N667, N5, N859);
nand NAND4 (N1863, N1859, N1745, N674, N1334);
buf BUF1 (N1864, N1862);
nand NAND4 (N1865, N1853, N149, N1501, N1799);
nor NOR3 (N1866, N1863, N1030, N1372);
nor NOR2 (N1867, N1864, N779);
xor XOR2 (N1868, N1857, N1069);
or OR3 (N1869, N1860, N1728, N578);
and AND4 (N1870, N1867, N728, N110, N217);
xor XOR2 (N1871, N1856, N1789);
buf BUF1 (N1872, N1869);
or OR3 (N1873, N1865, N363, N823);
xor XOR2 (N1874, N1861, N102);
buf BUF1 (N1875, N1839);
not NOT1 (N1876, N1868);
or OR3 (N1877, N1874, N1825, N245);
and AND4 (N1878, N1854, N349, N1850, N1572);
nand NAND2 (N1879, N1866, N763);
nand NAND2 (N1880, N1870, N265);
xor XOR2 (N1881, N1878, N939);
not NOT1 (N1882, N1871);
buf BUF1 (N1883, N1873);
nor NOR2 (N1884, N1881, N1863);
nor NOR3 (N1885, N1877, N1008, N659);
nand NAND2 (N1886, N1885, N1100);
nor NOR2 (N1887, N1886, N1860);
and AND3 (N1888, N1887, N1352, N491);
or OR3 (N1889, N1882, N1845, N844);
or OR4 (N1890, N1888, N554, N1793, N846);
not NOT1 (N1891, N1889);
buf BUF1 (N1892, N1880);
xor XOR2 (N1893, N1855, N1808);
nor NOR3 (N1894, N1872, N1727, N702);
nor NOR4 (N1895, N1893, N59, N613, N1177);
xor XOR2 (N1896, N1879, N1830);
and AND3 (N1897, N1876, N813, N1324);
xor XOR2 (N1898, N1894, N1594);
nand NAND3 (N1899, N1898, N1224, N183);
or OR3 (N1900, N1892, N377, N150);
or OR3 (N1901, N1883, N323, N1427);
nor NOR2 (N1902, N1884, N981);
nor NOR4 (N1903, N1896, N1600, N751, N1851);
buf BUF1 (N1904, N1890);
not NOT1 (N1905, N1903);
buf BUF1 (N1906, N1891);
buf BUF1 (N1907, N1901);
not NOT1 (N1908, N1895);
nor NOR4 (N1909, N1904, N1377, N1470, N1604);
not NOT1 (N1910, N1906);
nor NOR4 (N1911, N1902, N983, N1831, N257);
and AND4 (N1912, N1907, N1462, N1243, N451);
xor XOR2 (N1913, N1900, N232);
xor XOR2 (N1914, N1899, N1620);
not NOT1 (N1915, N1897);
buf BUF1 (N1916, N1912);
buf BUF1 (N1917, N1909);
buf BUF1 (N1918, N1910);
and AND4 (N1919, N1875, N1900, N479, N961);
or OR2 (N1920, N1918, N911);
nor NOR2 (N1921, N1917, N1594);
buf BUF1 (N1922, N1914);
or OR2 (N1923, N1922, N235);
xor XOR2 (N1924, N1915, N1709);
nor NOR2 (N1925, N1919, N1394);
nand NAND3 (N1926, N1913, N585, N446);
buf BUF1 (N1927, N1905);
not NOT1 (N1928, N1927);
nand NAND2 (N1929, N1908, N1817);
buf BUF1 (N1930, N1921);
xor XOR2 (N1931, N1923, N532);
nor NOR3 (N1932, N1920, N1000, N1192);
nor NOR4 (N1933, N1925, N32, N1114, N809);
nor NOR4 (N1934, N1911, N236, N774, N14);
buf BUF1 (N1935, N1934);
not NOT1 (N1936, N1928);
xor XOR2 (N1937, N1916, N92);
and AND2 (N1938, N1937, N1410);
nand NAND2 (N1939, N1935, N235);
buf BUF1 (N1940, N1932);
buf BUF1 (N1941, N1933);
not NOT1 (N1942, N1939);
buf BUF1 (N1943, N1929);
nand NAND3 (N1944, N1926, N486, N1922);
and AND3 (N1945, N1944, N41, N424);
or OR3 (N1946, N1940, N417, N457);
or OR2 (N1947, N1946, N1693);
buf BUF1 (N1948, N1938);
not NOT1 (N1949, N1930);
not NOT1 (N1950, N1941);
not NOT1 (N1951, N1945);
buf BUF1 (N1952, N1924);
not NOT1 (N1953, N1948);
nor NOR2 (N1954, N1931, N1027);
buf BUF1 (N1955, N1951);
nor NOR3 (N1956, N1955, N1890, N516);
and AND4 (N1957, N1949, N538, N1861, N1414);
buf BUF1 (N1958, N1950);
nand NAND3 (N1959, N1952, N16, N1428);
xor XOR2 (N1960, N1942, N1008);
and AND4 (N1961, N1959, N959, N1367, N1936);
xor XOR2 (N1962, N562, N1577);
xor XOR2 (N1963, N1954, N800);
and AND3 (N1964, N1957, N374, N1252);
buf BUF1 (N1965, N1962);
nor NOR3 (N1966, N1963, N497, N695);
or OR3 (N1967, N1960, N482, N806);
nor NOR2 (N1968, N1953, N1232);
xor XOR2 (N1969, N1943, N148);
and AND2 (N1970, N1967, N95);
or OR3 (N1971, N1968, N1240, N1961);
or OR2 (N1972, N1133, N1536);
not NOT1 (N1973, N1965);
not NOT1 (N1974, N1956);
or OR2 (N1975, N1972, N694);
nand NAND2 (N1976, N1969, N277);
or OR3 (N1977, N1973, N1819, N765);
and AND2 (N1978, N1958, N1430);
xor XOR2 (N1979, N1966, N415);
buf BUF1 (N1980, N1970);
buf BUF1 (N1981, N1978);
buf BUF1 (N1982, N1976);
nor NOR4 (N1983, N1964, N1157, N1712, N1406);
or OR2 (N1984, N1975, N544);
nor NOR2 (N1985, N1971, N1339);
and AND3 (N1986, N1985, N1479, N980);
and AND4 (N1987, N1986, N1245, N1222, N1860);
nand NAND3 (N1988, N1987, N1797, N83);
nand NAND4 (N1989, N1988, N1486, N271, N1846);
not NOT1 (N1990, N1979);
xor XOR2 (N1991, N1982, N550);
or OR3 (N1992, N1980, N710, N103);
buf BUF1 (N1993, N1983);
and AND2 (N1994, N1989, N980);
or OR4 (N1995, N1984, N1924, N801, N930);
or OR2 (N1996, N1974, N391);
xor XOR2 (N1997, N1994, N1224);
nand NAND2 (N1998, N1992, N54);
buf BUF1 (N1999, N1991);
not NOT1 (N2000, N1998);
and AND2 (N2001, N1977, N9);
nand NAND4 (N2002, N1996, N366, N385, N658);
nand NAND2 (N2003, N1995, N1665);
not NOT1 (N2004, N2001);
nand NAND3 (N2005, N2002, N597, N1010);
not NOT1 (N2006, N2005);
nand NAND4 (N2007, N2000, N192, N1234, N1370);
nor NOR4 (N2008, N2003, N1644, N639, N1007);
or OR4 (N2009, N1999, N743, N292, N1558);
nor NOR2 (N2010, N1990, N1440);
or OR3 (N2011, N1993, N1460, N892);
nor NOR4 (N2012, N2009, N931, N1578, N47);
nand NAND2 (N2013, N2008, N1360);
not NOT1 (N2014, N2012);
buf BUF1 (N2015, N2014);
nand NAND2 (N2016, N2013, N537);
xor XOR2 (N2017, N2016, N1467);
buf BUF1 (N2018, N2007);
xor XOR2 (N2019, N1947, N1651);
and AND4 (N2020, N2019, N1645, N1394, N212);
or OR3 (N2021, N2010, N1391, N1170);
or OR3 (N2022, N2006, N1716, N1279);
buf BUF1 (N2023, N1981);
or OR2 (N2024, N2004, N1730);
buf BUF1 (N2025, N2017);
buf BUF1 (N2026, N2023);
or OR3 (N2027, N2018, N1143, N764);
or OR3 (N2028, N2027, N1944, N2);
buf BUF1 (N2029, N2024);
or OR2 (N2030, N2028, N1078);
nand NAND4 (N2031, N1997, N1749, N571, N1938);
and AND3 (N2032, N2025, N721, N1806);
and AND4 (N2033, N2011, N1083, N1907, N546);
nor NOR3 (N2034, N2026, N1838, N688);
buf BUF1 (N2035, N2022);
not NOT1 (N2036, N2031);
nor NOR3 (N2037, N2021, N866, N618);
xor XOR2 (N2038, N2037, N361);
not NOT1 (N2039, N2033);
and AND2 (N2040, N2029, N711);
buf BUF1 (N2041, N2034);
xor XOR2 (N2042, N2040, N492);
nand NAND3 (N2043, N2032, N982, N1919);
or OR3 (N2044, N2038, N441, N537);
or OR3 (N2045, N2041, N435, N344);
nand NAND4 (N2046, N2043, N1403, N51, N1213);
nor NOR2 (N2047, N2036, N904);
nand NAND4 (N2048, N2039, N107, N1543, N1062);
not NOT1 (N2049, N2035);
buf BUF1 (N2050, N2049);
xor XOR2 (N2051, N2045, N1703);
nor NOR4 (N2052, N2044, N480, N1662, N568);
nand NAND4 (N2053, N2050, N1557, N942, N1874);
not NOT1 (N2054, N2015);
buf BUF1 (N2055, N2053);
buf BUF1 (N2056, N2054);
and AND4 (N2057, N2052, N1640, N1668, N762);
and AND3 (N2058, N2048, N1596, N160);
buf BUF1 (N2059, N2046);
nand NAND3 (N2060, N2042, N1626, N644);
and AND4 (N2061, N2047, N1983, N1262, N418);
buf BUF1 (N2062, N2058);
nand NAND4 (N2063, N2057, N336, N949, N1485);
buf BUF1 (N2064, N2062);
xor XOR2 (N2065, N2056, N1391);
or OR3 (N2066, N2020, N1070, N1869);
xor XOR2 (N2067, N2051, N1804);
not NOT1 (N2068, N2064);
not NOT1 (N2069, N2067);
and AND3 (N2070, N2055, N1641, N1287);
or OR3 (N2071, N2069, N1943, N540);
and AND2 (N2072, N2063, N407);
or OR3 (N2073, N2068, N1366, N1922);
and AND3 (N2074, N2065, N1535, N1857);
nor NOR3 (N2075, N2060, N1206, N498);
nand NAND4 (N2076, N2074, N1242, N26, N1431);
xor XOR2 (N2077, N2075, N778);
buf BUF1 (N2078, N2071);
not NOT1 (N2079, N2077);
and AND4 (N2080, N2066, N745, N1595, N875);
and AND2 (N2081, N2030, N1388);
or OR3 (N2082, N2073, N921, N446);
xor XOR2 (N2083, N2072, N1628);
not NOT1 (N2084, N2061);
and AND4 (N2085, N2059, N1162, N1271, N1795);
nor NOR3 (N2086, N2085, N675, N2016);
or OR3 (N2087, N2079, N982, N1805);
nand NAND4 (N2088, N2082, N1052, N214, N1950);
nor NOR2 (N2089, N2080, N1753);
or OR3 (N2090, N2086, N593, N1051);
nor NOR4 (N2091, N2090, N156, N26, N1669);
not NOT1 (N2092, N2070);
not NOT1 (N2093, N2089);
or OR4 (N2094, N2087, N1640, N859, N1055);
not NOT1 (N2095, N2076);
buf BUF1 (N2096, N2095);
or OR2 (N2097, N2092, N856);
nand NAND3 (N2098, N2091, N35, N1799);
xor XOR2 (N2099, N2097, N1131);
and AND4 (N2100, N2084, N1059, N1770, N1169);
nand NAND4 (N2101, N2099, N1137, N1171, N489);
not NOT1 (N2102, N2081);
nand NAND2 (N2103, N2102, N905);
or OR4 (N2104, N2088, N381, N576, N473);
xor XOR2 (N2105, N2083, N1329);
not NOT1 (N2106, N2094);
xor XOR2 (N2107, N2100, N1366);
and AND4 (N2108, N2096, N107, N927, N894);
not NOT1 (N2109, N2098);
nor NOR3 (N2110, N2108, N421, N1588);
nor NOR3 (N2111, N2106, N1283, N237);
nor NOR4 (N2112, N2110, N1725, N582, N529);
nand NAND3 (N2113, N2111, N1384, N356);
xor XOR2 (N2114, N2112, N1363);
xor XOR2 (N2115, N2103, N153);
and AND2 (N2116, N2115, N840);
or OR2 (N2117, N2104, N194);
or OR2 (N2118, N2101, N2045);
nand NAND4 (N2119, N2105, N948, N775, N1982);
or OR3 (N2120, N2117, N494, N1642);
nor NOR4 (N2121, N2118, N1958, N2063, N527);
nor NOR3 (N2122, N2107, N801, N1865);
and AND4 (N2123, N2109, N1470, N207, N1996);
buf BUF1 (N2124, N2113);
buf BUF1 (N2125, N2121);
or OR2 (N2126, N2122, N883);
and AND3 (N2127, N2116, N1961, N78);
xor XOR2 (N2128, N2093, N2100);
nand NAND3 (N2129, N2123, N1523, N480);
buf BUF1 (N2130, N2126);
nor NOR4 (N2131, N2127, N1967, N1923, N1743);
and AND4 (N2132, N2120, N651, N1824, N1819);
xor XOR2 (N2133, N2114, N958);
xor XOR2 (N2134, N2124, N2003);
nand NAND2 (N2135, N2130, N965);
and AND4 (N2136, N2131, N749, N624, N527);
nand NAND4 (N2137, N2129, N1189, N1669, N1596);
and AND4 (N2138, N2135, N716, N417, N1473);
buf BUF1 (N2139, N2137);
nand NAND4 (N2140, N2136, N97, N1217, N825);
nand NAND4 (N2141, N2078, N1217, N1910, N1953);
nor NOR4 (N2142, N2133, N803, N1758, N555);
or OR4 (N2143, N2138, N1083, N1586, N1089);
buf BUF1 (N2144, N2139);
buf BUF1 (N2145, N2143);
and AND4 (N2146, N2142, N969, N1792, N964);
xor XOR2 (N2147, N2145, N540);
nand NAND3 (N2148, N2125, N1582, N1000);
xor XOR2 (N2149, N2146, N1177);
or OR2 (N2150, N2149, N761);
nor NOR4 (N2151, N2144, N1951, N798, N926);
nand NAND3 (N2152, N2151, N1257, N282);
nand NAND3 (N2153, N2147, N1476, N1578);
or OR4 (N2154, N2153, N207, N1644, N1662);
buf BUF1 (N2155, N2152);
nand NAND4 (N2156, N2148, N2020, N1879, N1792);
nand NAND3 (N2157, N2154, N78, N55);
nor NOR2 (N2158, N2150, N2142);
xor XOR2 (N2159, N2156, N1464);
or OR3 (N2160, N2140, N2091, N665);
xor XOR2 (N2161, N2157, N1852);
and AND2 (N2162, N2160, N1548);
nand NAND3 (N2163, N2132, N585, N1846);
buf BUF1 (N2164, N2119);
buf BUF1 (N2165, N2162);
xor XOR2 (N2166, N2163, N699);
buf BUF1 (N2167, N2141);
not NOT1 (N2168, N2165);
or OR2 (N2169, N2167, N722);
or OR2 (N2170, N2164, N978);
nor NOR2 (N2171, N2169, N286);
and AND3 (N2172, N2128, N1518, N2073);
not NOT1 (N2173, N2134);
nand NAND3 (N2174, N2159, N150, N891);
or OR4 (N2175, N2171, N921, N1402, N930);
nand NAND2 (N2176, N2168, N68);
buf BUF1 (N2177, N2161);
xor XOR2 (N2178, N2172, N800);
nand NAND4 (N2179, N2177, N1994, N1167, N1498);
xor XOR2 (N2180, N2170, N2029);
xor XOR2 (N2181, N2174, N444);
and AND3 (N2182, N2158, N966, N594);
buf BUF1 (N2183, N2179);
xor XOR2 (N2184, N2173, N473);
and AND2 (N2185, N2181, N2126);
or OR4 (N2186, N2180, N261, N1649, N731);
xor XOR2 (N2187, N2176, N1516);
xor XOR2 (N2188, N2187, N1683);
and AND2 (N2189, N2166, N2031);
nand NAND2 (N2190, N2184, N1464);
not NOT1 (N2191, N2189);
or OR3 (N2192, N2191, N1925, N1567);
buf BUF1 (N2193, N2190);
nor NOR3 (N2194, N2175, N835, N12);
nor NOR3 (N2195, N2188, N1012, N188);
nand NAND4 (N2196, N2194, N434, N1688, N1893);
nand NAND4 (N2197, N2183, N265, N1819, N2174);
nor NOR4 (N2198, N2192, N869, N1133, N885);
and AND2 (N2199, N2155, N36);
and AND4 (N2200, N2199, N2198, N1706, N1072);
buf BUF1 (N2201, N1945);
or OR2 (N2202, N2178, N1898);
and AND4 (N2203, N2186, N1686, N1564, N1371);
not NOT1 (N2204, N2197);
xor XOR2 (N2205, N2195, N105);
nand NAND2 (N2206, N2203, N1199);
or OR4 (N2207, N2206, N1267, N1818, N2151);
and AND3 (N2208, N2207, N460, N1539);
nand NAND2 (N2209, N2205, N43);
xor XOR2 (N2210, N2193, N234);
buf BUF1 (N2211, N2182);
and AND4 (N2212, N2200, N94, N801, N160);
and AND2 (N2213, N2196, N2199);
not NOT1 (N2214, N2185);
nor NOR2 (N2215, N2209, N1177);
or OR4 (N2216, N2204, N1418, N2039, N370);
and AND3 (N2217, N2210, N1664, N775);
or OR2 (N2218, N2216, N1372);
or OR2 (N2219, N2201, N134);
nand NAND3 (N2220, N2202, N2077, N852);
not NOT1 (N2221, N2208);
nand NAND2 (N2222, N2220, N519);
nand NAND4 (N2223, N2214, N113, N91, N1776);
and AND3 (N2224, N2217, N333, N1383);
and AND3 (N2225, N2222, N1439, N1);
xor XOR2 (N2226, N2223, N144);
or OR2 (N2227, N2212, N237);
not NOT1 (N2228, N2211);
not NOT1 (N2229, N2221);
not NOT1 (N2230, N2228);
xor XOR2 (N2231, N2226, N2008);
and AND4 (N2232, N2215, N1756, N805, N1716);
and AND2 (N2233, N2225, N1397);
or OR3 (N2234, N2227, N1637, N773);
and AND2 (N2235, N2232, N1927);
nor NOR3 (N2236, N2218, N583, N927);
xor XOR2 (N2237, N2231, N1303);
and AND2 (N2238, N2213, N1449);
or OR3 (N2239, N2238, N2000, N822);
not NOT1 (N2240, N2219);
and AND4 (N2241, N2237, N666, N517, N407);
buf BUF1 (N2242, N2241);
buf BUF1 (N2243, N2234);
xor XOR2 (N2244, N2236, N1892);
nand NAND4 (N2245, N2233, N1789, N108, N1210);
nor NOR4 (N2246, N2240, N550, N372, N1753);
nor NOR2 (N2247, N2239, N2131);
nand NAND3 (N2248, N2224, N703, N2236);
xor XOR2 (N2249, N2235, N1848);
nand NAND4 (N2250, N2230, N1935, N165, N1238);
buf BUF1 (N2251, N2243);
xor XOR2 (N2252, N2245, N63);
nor NOR3 (N2253, N2229, N2004, N910);
not NOT1 (N2254, N2253);
or OR3 (N2255, N2252, N730, N799);
nand NAND2 (N2256, N2251, N746);
xor XOR2 (N2257, N2242, N281);
nor NOR4 (N2258, N2247, N1025, N1193, N2184);
buf BUF1 (N2259, N2254);
buf BUF1 (N2260, N2250);
nand NAND4 (N2261, N2258, N54, N2177, N703);
nand NAND3 (N2262, N2259, N1544, N536);
nor NOR3 (N2263, N2249, N1376, N1936);
and AND4 (N2264, N2257, N1089, N800, N1557);
buf BUF1 (N2265, N2260);
xor XOR2 (N2266, N2255, N519);
and AND3 (N2267, N2262, N1544, N207);
buf BUF1 (N2268, N2264);
not NOT1 (N2269, N2248);
nor NOR4 (N2270, N2268, N1662, N1745, N1689);
or OR4 (N2271, N2263, N2079, N1952, N934);
nand NAND2 (N2272, N2246, N541);
nor NOR3 (N2273, N2265, N770, N13);
xor XOR2 (N2274, N2273, N296);
or OR2 (N2275, N2274, N1487);
buf BUF1 (N2276, N2271);
or OR3 (N2277, N2270, N922, N1814);
xor XOR2 (N2278, N2267, N885);
buf BUF1 (N2279, N2272);
or OR2 (N2280, N2261, N109);
nor NOR3 (N2281, N2276, N1496, N308);
buf BUF1 (N2282, N2278);
nor NOR4 (N2283, N2266, N34, N532, N1834);
xor XOR2 (N2284, N2269, N662);
and AND2 (N2285, N2279, N1779);
buf BUF1 (N2286, N2280);
nand NAND4 (N2287, N2277, N639, N1074, N334);
and AND4 (N2288, N2283, N22, N699, N1099);
buf BUF1 (N2289, N2256);
nor NOR3 (N2290, N2286, N1537, N1442);
nand NAND4 (N2291, N2287, N1658, N1592, N981);
buf BUF1 (N2292, N2291);
xor XOR2 (N2293, N2284, N142);
and AND3 (N2294, N2290, N515, N140);
and AND4 (N2295, N2289, N1813, N383, N1600);
buf BUF1 (N2296, N2295);
buf BUF1 (N2297, N2296);
or OR2 (N2298, N2244, N1981);
nor NOR4 (N2299, N2288, N2154, N1916, N2285);
nand NAND3 (N2300, N1909, N152, N2136);
not NOT1 (N2301, N2297);
nor NOR2 (N2302, N2300, N1709);
nand NAND4 (N2303, N2301, N176, N1450, N2081);
not NOT1 (N2304, N2281);
and AND4 (N2305, N2282, N298, N1543, N1594);
and AND3 (N2306, N2305, N74, N1768);
xor XOR2 (N2307, N2304, N1888);
nor NOR4 (N2308, N2292, N1505, N2066, N1561);
not NOT1 (N2309, N2298);
xor XOR2 (N2310, N2293, N383);
not NOT1 (N2311, N2294);
nand NAND4 (N2312, N2308, N883, N2108, N1707);
or OR4 (N2313, N2311, N568, N1718, N1523);
buf BUF1 (N2314, N2299);
buf BUF1 (N2315, N2303);
or OR4 (N2316, N2314, N1991, N423, N924);
or OR2 (N2317, N2309, N1517);
buf BUF1 (N2318, N2306);
and AND2 (N2319, N2307, N38);
not NOT1 (N2320, N2310);
nand NAND4 (N2321, N2316, N1012, N1673, N1137);
nand NAND3 (N2322, N2319, N993, N1868);
and AND3 (N2323, N2320, N1114, N2070);
xor XOR2 (N2324, N2312, N1367);
xor XOR2 (N2325, N2324, N2276);
and AND2 (N2326, N2318, N1168);
nor NOR4 (N2327, N2321, N1868, N1195, N1422);
not NOT1 (N2328, N2323);
or OR4 (N2329, N2313, N598, N2120, N1053);
and AND4 (N2330, N2275, N1974, N1662, N874);
nand NAND3 (N2331, N2326, N2281, N784);
not NOT1 (N2332, N2317);
not NOT1 (N2333, N2325);
buf BUF1 (N2334, N2328);
buf BUF1 (N2335, N2302);
and AND3 (N2336, N2329, N292, N1020);
buf BUF1 (N2337, N2322);
buf BUF1 (N2338, N2315);
buf BUF1 (N2339, N2335);
or OR4 (N2340, N2330, N2298, N35, N1189);
xor XOR2 (N2341, N2337, N450);
not NOT1 (N2342, N2341);
buf BUF1 (N2343, N2332);
buf BUF1 (N2344, N2340);
or OR3 (N2345, N2327, N1649, N2133);
nand NAND4 (N2346, N2336, N2345, N962, N146);
buf BUF1 (N2347, N747);
or OR2 (N2348, N2346, N2327);
buf BUF1 (N2349, N2347);
nor NOR3 (N2350, N2342, N1660, N1810);
nand NAND2 (N2351, N2339, N546);
xor XOR2 (N2352, N2344, N2341);
buf BUF1 (N2353, N2351);
nand NAND4 (N2354, N2352, N309, N6, N2059);
nand NAND2 (N2355, N2331, N612);
nand NAND3 (N2356, N2355, N2214, N1075);
buf BUF1 (N2357, N2338);
xor XOR2 (N2358, N2350, N2131);
and AND3 (N2359, N2356, N1937, N1990);
not NOT1 (N2360, N2359);
nor NOR4 (N2361, N2360, N1587, N1380, N4);
not NOT1 (N2362, N2353);
and AND2 (N2363, N2333, N50);
xor XOR2 (N2364, N2349, N1013);
or OR3 (N2365, N2357, N2324, N751);
xor XOR2 (N2366, N2361, N2216);
buf BUF1 (N2367, N2358);
nor NOR3 (N2368, N2343, N1643, N386);
not NOT1 (N2369, N2367);
buf BUF1 (N2370, N2334);
buf BUF1 (N2371, N2348);
or OR4 (N2372, N2366, N2330, N537, N1922);
buf BUF1 (N2373, N2372);
xor XOR2 (N2374, N2370, N1515);
buf BUF1 (N2375, N2368);
and AND2 (N2376, N2354, N2116);
nor NOR2 (N2377, N2362, N2160);
and AND2 (N2378, N2365, N1788);
nor NOR3 (N2379, N2369, N69, N237);
nand NAND3 (N2380, N2378, N1006, N318);
or OR4 (N2381, N2371, N1896, N1356, N296);
not NOT1 (N2382, N2376);
not NOT1 (N2383, N2363);
xor XOR2 (N2384, N2380, N627);
not NOT1 (N2385, N2375);
or OR2 (N2386, N2383, N389);
nand NAND3 (N2387, N2364, N819, N691);
nor NOR4 (N2388, N2377, N2156, N236, N487);
nor NOR2 (N2389, N2374, N1580);
nand NAND2 (N2390, N2388, N996);
buf BUF1 (N2391, N2384);
xor XOR2 (N2392, N2389, N804);
buf BUF1 (N2393, N2381);
not NOT1 (N2394, N2385);
or OR2 (N2395, N2379, N1870);
nor NOR2 (N2396, N2391, N1262);
xor XOR2 (N2397, N2382, N2052);
and AND3 (N2398, N2386, N65, N320);
xor XOR2 (N2399, N2392, N2070);
buf BUF1 (N2400, N2390);
xor XOR2 (N2401, N2394, N2105);
and AND3 (N2402, N2399, N1549, N2191);
not NOT1 (N2403, N2401);
nand NAND2 (N2404, N2393, N270);
buf BUF1 (N2405, N2400);
xor XOR2 (N2406, N2402, N93);
or OR4 (N2407, N2404, N762, N2275, N2375);
and AND2 (N2408, N2395, N1297);
not NOT1 (N2409, N2403);
not NOT1 (N2410, N2397);
not NOT1 (N2411, N2406);
nor NOR2 (N2412, N2405, N1434);
buf BUF1 (N2413, N2387);
or OR2 (N2414, N2407, N1220);
or OR2 (N2415, N2413, N1059);
and AND3 (N2416, N2415, N1527, N166);
and AND2 (N2417, N2409, N1527);
and AND4 (N2418, N2408, N1210, N2267, N359);
xor XOR2 (N2419, N2396, N996);
nand NAND2 (N2420, N2414, N1519);
xor XOR2 (N2421, N2410, N74);
nor NOR2 (N2422, N2373, N1670);
buf BUF1 (N2423, N2421);
and AND4 (N2424, N2417, N1503, N148, N1056);
not NOT1 (N2425, N2418);
and AND4 (N2426, N2425, N1369, N123, N2112);
nand NAND2 (N2427, N2411, N928);
nor NOR4 (N2428, N2416, N1970, N370, N989);
or OR3 (N2429, N2398, N1403, N1276);
buf BUF1 (N2430, N2429);
xor XOR2 (N2431, N2422, N1675);
or OR4 (N2432, N2431, N1865, N1062, N803);
xor XOR2 (N2433, N2423, N981);
nor NOR2 (N2434, N2424, N2373);
not NOT1 (N2435, N2428);
or OR2 (N2436, N2433, N650);
nor NOR4 (N2437, N2436, N2210, N1883, N2060);
nand NAND4 (N2438, N2435, N1880, N1546, N534);
xor XOR2 (N2439, N2420, N1629);
nor NOR2 (N2440, N2439, N63);
xor XOR2 (N2441, N2427, N2280);
buf BUF1 (N2442, N2430);
or OR2 (N2443, N2440, N958);
nor NOR3 (N2444, N2443, N2084, N165);
nand NAND4 (N2445, N2442, N307, N35, N1882);
nand NAND3 (N2446, N2426, N1518, N920);
or OR4 (N2447, N2437, N2366, N526, N1867);
and AND4 (N2448, N2446, N740, N1214, N458);
nand NAND4 (N2449, N2444, N1720, N1618, N201);
not NOT1 (N2450, N2434);
nand NAND2 (N2451, N2445, N748);
nor NOR4 (N2452, N2419, N2072, N2036, N1826);
not NOT1 (N2453, N2441);
and AND4 (N2454, N2432, N114, N1694, N1398);
xor XOR2 (N2455, N2448, N1228);
nand NAND4 (N2456, N2452, N2176, N2144, N1643);
not NOT1 (N2457, N2454);
and AND2 (N2458, N2453, N590);
nand NAND2 (N2459, N2412, N1799);
nor NOR2 (N2460, N2456, N348);
and AND3 (N2461, N2449, N1569, N488);
or OR4 (N2462, N2459, N224, N678, N1512);
and AND4 (N2463, N2451, N471, N1465, N1086);
not NOT1 (N2464, N2461);
buf BUF1 (N2465, N2458);
xor XOR2 (N2466, N2464, N488);
or OR4 (N2467, N2462, N1495, N1174, N1262);
xor XOR2 (N2468, N2438, N1729);
and AND4 (N2469, N2467, N106, N553, N2092);
nand NAND2 (N2470, N2465, N1275);
xor XOR2 (N2471, N2470, N2378);
and AND2 (N2472, N2457, N2187);
not NOT1 (N2473, N2463);
or OR4 (N2474, N2469, N846, N2242, N871);
or OR2 (N2475, N2474, N894);
nand NAND4 (N2476, N2447, N736, N479, N2166);
xor XOR2 (N2477, N2473, N2162);
and AND3 (N2478, N2471, N1155, N1440);
or OR2 (N2479, N2478, N2469);
or OR4 (N2480, N2477, N1040, N457, N284);
not NOT1 (N2481, N2476);
and AND3 (N2482, N2472, N2163, N1079);
xor XOR2 (N2483, N2450, N1318);
buf BUF1 (N2484, N2481);
not NOT1 (N2485, N2484);
or OR2 (N2486, N2482, N2296);
not NOT1 (N2487, N2480);
nor NOR2 (N2488, N2485, N1935);
nor NOR4 (N2489, N2475, N393, N1618, N182);
nor NOR3 (N2490, N2479, N1040, N2251);
and AND2 (N2491, N2490, N1493);
buf BUF1 (N2492, N2455);
nor NOR3 (N2493, N2483, N689, N982);
nand NAND4 (N2494, N2489, N642, N1231, N28);
nand NAND2 (N2495, N2460, N2254);
nand NAND2 (N2496, N2488, N1160);
and AND2 (N2497, N2494, N30);
or OR2 (N2498, N2497, N140);
nand NAND4 (N2499, N2498, N1576, N1029, N39);
not NOT1 (N2500, N2496);
buf BUF1 (N2501, N2468);
and AND2 (N2502, N2491, N607);
not NOT1 (N2503, N2500);
xor XOR2 (N2504, N2501, N2173);
or OR3 (N2505, N2499, N655, N1074);
and AND4 (N2506, N2493, N2314, N1378, N1855);
or OR3 (N2507, N2487, N22, N1588);
buf BUF1 (N2508, N2507);
and AND3 (N2509, N2466, N1986, N146);
nand NAND3 (N2510, N2486, N1617, N2281);
xor XOR2 (N2511, N2508, N1389);
nand NAND3 (N2512, N2502, N1433, N1939);
not NOT1 (N2513, N2504);
buf BUF1 (N2514, N2503);
buf BUF1 (N2515, N2492);
nor NOR3 (N2516, N2513, N2382, N1731);
and AND3 (N2517, N2495, N1535, N1225);
nand NAND4 (N2518, N2517, N1647, N2275, N1525);
xor XOR2 (N2519, N2510, N2022);
not NOT1 (N2520, N2505);
and AND4 (N2521, N2519, N753, N830, N1087);
nand NAND3 (N2522, N2514, N1519, N36);
not NOT1 (N2523, N2509);
and AND3 (N2524, N2521, N1826, N10);
nor NOR2 (N2525, N2520, N876);
nor NOR4 (N2526, N2523, N698, N911, N2263);
buf BUF1 (N2527, N2525);
nand NAND3 (N2528, N2506, N245, N2459);
nand NAND3 (N2529, N2522, N1603, N902);
nand NAND4 (N2530, N2529, N214, N2238, N151);
xor XOR2 (N2531, N2526, N1016);
nor NOR3 (N2532, N2531, N1682, N1437);
xor XOR2 (N2533, N2527, N443);
or OR4 (N2534, N2516, N1902, N1593, N7);
nand NAND3 (N2535, N2512, N311, N933);
not NOT1 (N2536, N2524);
not NOT1 (N2537, N2511);
or OR2 (N2538, N2515, N991);
xor XOR2 (N2539, N2532, N2342);
nor NOR3 (N2540, N2534, N1479, N2252);
nand NAND4 (N2541, N2539, N1429, N1783, N205);
not NOT1 (N2542, N2538);
nand NAND2 (N2543, N2518, N1669);
nor NOR4 (N2544, N2533, N673, N1806, N1965);
nor NOR2 (N2545, N2541, N1371);
nand NAND4 (N2546, N2543, N1983, N1534, N777);
buf BUF1 (N2547, N2536);
nand NAND4 (N2548, N2540, N1614, N1954, N1996);
nand NAND2 (N2549, N2542, N1653);
and AND4 (N2550, N2546, N100, N2409, N551);
and AND4 (N2551, N2548, N1567, N1434, N341);
xor XOR2 (N2552, N2549, N2201);
nor NOR2 (N2553, N2545, N1439);
buf BUF1 (N2554, N2547);
nand NAND2 (N2555, N2551, N572);
and AND2 (N2556, N2537, N553);
nor NOR2 (N2557, N2550, N651);
nand NAND4 (N2558, N2552, N1541, N2259, N1418);
xor XOR2 (N2559, N2530, N1946);
or OR2 (N2560, N2528, N780);
nor NOR4 (N2561, N2556, N1629, N978, N454);
and AND4 (N2562, N2559, N1507, N2072, N2134);
or OR2 (N2563, N2553, N533);
and AND3 (N2564, N2544, N1241, N1111);
buf BUF1 (N2565, N2564);
xor XOR2 (N2566, N2535, N1155);
buf BUF1 (N2567, N2557);
or OR3 (N2568, N2566, N1748, N1353);
xor XOR2 (N2569, N2558, N389);
not NOT1 (N2570, N2560);
buf BUF1 (N2571, N2570);
or OR2 (N2572, N2571, N547);
and AND2 (N2573, N2555, N1288);
or OR2 (N2574, N2563, N1710);
nand NAND2 (N2575, N2572, N413);
xor XOR2 (N2576, N2561, N2441);
nor NOR3 (N2577, N2575, N2400, N1369);
buf BUF1 (N2578, N2573);
buf BUF1 (N2579, N2569);
nor NOR2 (N2580, N2574, N1537);
or OR2 (N2581, N2579, N18);
or OR4 (N2582, N2554, N1972, N1658, N2111);
and AND2 (N2583, N2568, N1855);
or OR4 (N2584, N2562, N992, N1778, N56);
xor XOR2 (N2585, N2582, N1270);
or OR3 (N2586, N2576, N1640, N1638);
nand NAND4 (N2587, N2578, N2372, N1083, N1757);
or OR4 (N2588, N2586, N693, N2443, N417);
not NOT1 (N2589, N2581);
not NOT1 (N2590, N2584);
nor NOR2 (N2591, N2585, N503);
buf BUF1 (N2592, N2565);
nor NOR4 (N2593, N2580, N775, N373, N621);
not NOT1 (N2594, N2589);
or OR3 (N2595, N2592, N767, N2384);
nor NOR4 (N2596, N2591, N2584, N2217, N118);
or OR4 (N2597, N2590, N897, N2109, N1357);
nor NOR4 (N2598, N2587, N1787, N474, N810);
buf BUF1 (N2599, N2598);
xor XOR2 (N2600, N2588, N443);
and AND2 (N2601, N2597, N335);
not NOT1 (N2602, N2583);
not NOT1 (N2603, N2596);
nand NAND3 (N2604, N2593, N264, N475);
buf BUF1 (N2605, N2602);
and AND3 (N2606, N2603, N753, N1875);
and AND2 (N2607, N2577, N817);
and AND2 (N2608, N2595, N480);
nor NOR3 (N2609, N2601, N658, N1573);
and AND2 (N2610, N2605, N9);
xor XOR2 (N2611, N2607, N2249);
or OR2 (N2612, N2594, N438);
and AND2 (N2613, N2612, N1019);
xor XOR2 (N2614, N2613, N2329);
nor NOR3 (N2615, N2599, N1643, N2008);
buf BUF1 (N2616, N2611);
nand NAND3 (N2617, N2610, N2356, N436);
or OR2 (N2618, N2614, N1147);
nor NOR3 (N2619, N2615, N1547, N2482);
xor XOR2 (N2620, N2567, N1730);
nor NOR2 (N2621, N2608, N835);
nand NAND3 (N2622, N2619, N1693, N1653);
buf BUF1 (N2623, N2620);
or OR3 (N2624, N2623, N1837, N1832);
and AND4 (N2625, N2622, N956, N1927, N1516);
not NOT1 (N2626, N2617);
and AND3 (N2627, N2624, N671, N2623);
or OR4 (N2628, N2600, N1013, N2007, N488);
not NOT1 (N2629, N2628);
nand NAND4 (N2630, N2604, N2475, N686, N1091);
and AND2 (N2631, N2626, N2156);
nor NOR3 (N2632, N2606, N1692, N1573);
xor XOR2 (N2633, N2616, N1116);
or OR3 (N2634, N2621, N1161, N3);
nor NOR2 (N2635, N2618, N230);
nor NOR3 (N2636, N2630, N2364, N2159);
nor NOR3 (N2637, N2609, N317, N1784);
or OR3 (N2638, N2632, N486, N797);
or OR4 (N2639, N2637, N2009, N1204, N1817);
or OR2 (N2640, N2635, N696);
buf BUF1 (N2641, N2639);
buf BUF1 (N2642, N2625);
not NOT1 (N2643, N2631);
and AND2 (N2644, N2633, N2544);
not NOT1 (N2645, N2641);
and AND2 (N2646, N2640, N2324);
and AND4 (N2647, N2643, N211, N816, N283);
buf BUF1 (N2648, N2646);
and AND4 (N2649, N2638, N1352, N619, N702);
and AND2 (N2650, N2627, N2004);
nor NOR4 (N2651, N2647, N984, N834, N2582);
nand NAND2 (N2652, N2651, N1820);
xor XOR2 (N2653, N2648, N2061);
nand NAND2 (N2654, N2652, N1023);
nor NOR2 (N2655, N2654, N1552);
buf BUF1 (N2656, N2634);
not NOT1 (N2657, N2653);
and AND4 (N2658, N2636, N707, N1116, N1132);
xor XOR2 (N2659, N2657, N974);
nand NAND3 (N2660, N2642, N650, N259);
and AND3 (N2661, N2644, N2035, N544);
buf BUF1 (N2662, N2655);
nor NOR2 (N2663, N2656, N1780);
not NOT1 (N2664, N2662);
buf BUF1 (N2665, N2650);
xor XOR2 (N2666, N2660, N1313);
xor XOR2 (N2667, N2645, N719);
nand NAND2 (N2668, N2659, N1303);
not NOT1 (N2669, N2665);
nor NOR3 (N2670, N2658, N2179, N782);
nor NOR2 (N2671, N2670, N8);
not NOT1 (N2672, N2668);
buf BUF1 (N2673, N2629);
nor NOR4 (N2674, N2661, N816, N920, N1578);
nor NOR4 (N2675, N2664, N2427, N1948, N127);
buf BUF1 (N2676, N2666);
nor NOR4 (N2677, N2672, N665, N2636, N1254);
nor NOR2 (N2678, N2677, N2450);
and AND4 (N2679, N2671, N2524, N1596, N74);
xor XOR2 (N2680, N2678, N2223);
or OR3 (N2681, N2667, N2401, N1957);
buf BUF1 (N2682, N2675);
nor NOR3 (N2683, N2673, N486, N1822);
and AND3 (N2684, N2676, N2526, N2285);
buf BUF1 (N2685, N2669);
not NOT1 (N2686, N2649);
or OR3 (N2687, N2663, N2471, N477);
and AND3 (N2688, N2682, N125, N1164);
and AND3 (N2689, N2687, N246, N20);
not NOT1 (N2690, N2680);
or OR3 (N2691, N2688, N1656, N2400);
or OR3 (N2692, N2691, N1671, N2229);
not NOT1 (N2693, N2689);
nand NAND4 (N2694, N2685, N2025, N497, N2450);
and AND2 (N2695, N2694, N105);
nor NOR4 (N2696, N2684, N1546, N1456, N480);
buf BUF1 (N2697, N2693);
and AND2 (N2698, N2679, N417);
xor XOR2 (N2699, N2692, N1836);
or OR2 (N2700, N2683, N1395);
or OR3 (N2701, N2690, N162, N381);
nand NAND3 (N2702, N2700, N2466, N2365);
not NOT1 (N2703, N2696);
and AND4 (N2704, N2695, N2696, N2315, N1845);
buf BUF1 (N2705, N2686);
nand NAND2 (N2706, N2702, N532);
buf BUF1 (N2707, N2701);
nand NAND2 (N2708, N2699, N2486);
not NOT1 (N2709, N2706);
not NOT1 (N2710, N2707);
nand NAND3 (N2711, N2698, N1128, N2070);
nand NAND3 (N2712, N2704, N1166, N1967);
not NOT1 (N2713, N2711);
nor NOR3 (N2714, N2712, N2643, N1937);
buf BUF1 (N2715, N2705);
nor NOR2 (N2716, N2674, N2605);
xor XOR2 (N2717, N2710, N1);
or OR2 (N2718, N2697, N1258);
not NOT1 (N2719, N2716);
xor XOR2 (N2720, N2708, N2304);
not NOT1 (N2721, N2709);
and AND3 (N2722, N2721, N1465, N408);
nand NAND4 (N2723, N2681, N542, N882, N2218);
nor NOR4 (N2724, N2703, N955, N655, N962);
nor NOR4 (N2725, N2715, N1222, N1304, N1616);
buf BUF1 (N2726, N2714);
nor NOR4 (N2727, N2717, N2087, N693, N572);
xor XOR2 (N2728, N2713, N2612);
nand NAND3 (N2729, N2723, N625, N31);
or OR3 (N2730, N2725, N355, N1426);
xor XOR2 (N2731, N2727, N2634);
xor XOR2 (N2732, N2724, N972);
and AND2 (N2733, N2729, N2053);
and AND4 (N2734, N2730, N2141, N2636, N2548);
not NOT1 (N2735, N2720);
xor XOR2 (N2736, N2731, N865);
not NOT1 (N2737, N2728);
nand NAND4 (N2738, N2726, N222, N1120, N2235);
xor XOR2 (N2739, N2734, N721);
xor XOR2 (N2740, N2719, N26);
nor NOR3 (N2741, N2740, N882, N234);
and AND3 (N2742, N2741, N234, N14);
and AND3 (N2743, N2732, N954, N4);
not NOT1 (N2744, N2735);
or OR2 (N2745, N2738, N502);
not NOT1 (N2746, N2733);
and AND2 (N2747, N2722, N762);
xor XOR2 (N2748, N2736, N223);
xor XOR2 (N2749, N2718, N624);
or OR4 (N2750, N2746, N2030, N161, N977);
nor NOR4 (N2751, N2737, N882, N2351, N1323);
not NOT1 (N2752, N2750);
or OR3 (N2753, N2751, N90, N623);
nor NOR4 (N2754, N2747, N2699, N2277, N2252);
xor XOR2 (N2755, N2749, N925);
not NOT1 (N2756, N2752);
nand NAND2 (N2757, N2742, N1104);
nand NAND2 (N2758, N2755, N160);
not NOT1 (N2759, N2745);
or OR2 (N2760, N2744, N236);
not NOT1 (N2761, N2753);
buf BUF1 (N2762, N2754);
xor XOR2 (N2763, N2743, N1980);
or OR2 (N2764, N2759, N802);
nand NAND4 (N2765, N2763, N2730, N2204, N1103);
xor XOR2 (N2766, N2764, N2097);
nand NAND3 (N2767, N2760, N1170, N2322);
not NOT1 (N2768, N2761);
nand NAND3 (N2769, N2766, N2075, N544);
buf BUF1 (N2770, N2758);
nor NOR4 (N2771, N2756, N746, N2156, N95);
or OR2 (N2772, N2757, N443);
buf BUF1 (N2773, N2739);
buf BUF1 (N2774, N2773);
not NOT1 (N2775, N2769);
nand NAND4 (N2776, N2765, N291, N1834, N1249);
or OR2 (N2777, N2774, N658);
and AND2 (N2778, N2776, N1711);
not NOT1 (N2779, N2778);
nor NOR2 (N2780, N2777, N2513);
and AND4 (N2781, N2779, N2504, N2295, N2678);
nor NOR4 (N2782, N2771, N758, N1416, N1631);
buf BUF1 (N2783, N2762);
nand NAND2 (N2784, N2768, N2026);
nor NOR4 (N2785, N2784, N526, N12, N2378);
not NOT1 (N2786, N2772);
and AND4 (N2787, N2782, N1979, N1910, N813);
not NOT1 (N2788, N2786);
not NOT1 (N2789, N2767);
nand NAND3 (N2790, N2787, N1343, N2667);
nor NOR3 (N2791, N2780, N2771, N1193);
nand NAND4 (N2792, N2783, N2492, N1480, N1562);
xor XOR2 (N2793, N2785, N1532);
nor NOR2 (N2794, N2788, N1450);
nand NAND3 (N2795, N2790, N2728, N2305);
and AND3 (N2796, N2793, N1685, N266);
nor NOR3 (N2797, N2781, N1820, N709);
nand NAND3 (N2798, N2789, N1720, N2239);
buf BUF1 (N2799, N2791);
nor NOR3 (N2800, N2794, N538, N2101);
xor XOR2 (N2801, N2770, N2066);
or OR2 (N2802, N2795, N1954);
or OR3 (N2803, N2792, N787, N2633);
buf BUF1 (N2804, N2803);
or OR3 (N2805, N2748, N929, N2787);
not NOT1 (N2806, N2797);
nand NAND2 (N2807, N2800, N2448);
and AND2 (N2808, N2775, N1563);
buf BUF1 (N2809, N2798);
nor NOR3 (N2810, N2806, N666, N1785);
or OR3 (N2811, N2807, N698, N805);
xor XOR2 (N2812, N2802, N2130);
not NOT1 (N2813, N2799);
and AND4 (N2814, N2808, N2125, N1752, N2034);
and AND2 (N2815, N2810, N906);
and AND4 (N2816, N2805, N920, N31, N1208);
or OR3 (N2817, N2811, N610, N1360);
not NOT1 (N2818, N2801);
or OR3 (N2819, N2796, N456, N1362);
xor XOR2 (N2820, N2814, N773);
and AND3 (N2821, N2812, N956, N1570);
buf BUF1 (N2822, N2817);
nor NOR3 (N2823, N2816, N608, N2187);
or OR2 (N2824, N2809, N332);
xor XOR2 (N2825, N2824, N907);
xor XOR2 (N2826, N2815, N2319);
not NOT1 (N2827, N2820);
and AND2 (N2828, N2804, N1394);
and AND4 (N2829, N2813, N613, N2293, N181);
xor XOR2 (N2830, N2826, N2414);
or OR2 (N2831, N2819, N1906);
not NOT1 (N2832, N2828);
nand NAND3 (N2833, N2831, N276, N178);
buf BUF1 (N2834, N2823);
xor XOR2 (N2835, N2834, N2261);
xor XOR2 (N2836, N2835, N838);
and AND3 (N2837, N2822, N2474, N2058);
nand NAND2 (N2838, N2825, N2812);
and AND4 (N2839, N2833, N1402, N1859, N633);
not NOT1 (N2840, N2837);
nor NOR4 (N2841, N2830, N2383, N479, N421);
nand NAND3 (N2842, N2827, N2268, N759);
not NOT1 (N2843, N2829);
and AND4 (N2844, N2821, N331, N63, N211);
nor NOR4 (N2845, N2832, N2060, N1257, N409);
nor NOR4 (N2846, N2841, N356, N2845, N899);
and AND2 (N2847, N1971, N2216);
not NOT1 (N2848, N2842);
nand NAND3 (N2849, N2839, N903, N1367);
xor XOR2 (N2850, N2838, N2497);
buf BUF1 (N2851, N2843);
xor XOR2 (N2852, N2848, N401);
and AND3 (N2853, N2850, N1698, N387);
xor XOR2 (N2854, N2818, N2732);
nand NAND3 (N2855, N2852, N1997, N1119);
or OR4 (N2856, N2854, N334, N840, N2693);
and AND4 (N2857, N2855, N1264, N1891, N548);
nor NOR3 (N2858, N2857, N2200, N2630);
not NOT1 (N2859, N2858);
not NOT1 (N2860, N2847);
buf BUF1 (N2861, N2851);
not NOT1 (N2862, N2840);
xor XOR2 (N2863, N2859, N2791);
and AND2 (N2864, N2836, N2149);
nand NAND2 (N2865, N2862, N2696);
buf BUF1 (N2866, N2853);
or OR3 (N2867, N2863, N1690, N731);
or OR4 (N2868, N2866, N71, N2062, N2843);
xor XOR2 (N2869, N2864, N513);
nand NAND2 (N2870, N2856, N1356);
not NOT1 (N2871, N2869);
or OR4 (N2872, N2868, N147, N1003, N1651);
nand NAND2 (N2873, N2861, N2098);
xor XOR2 (N2874, N2870, N1402);
nand NAND3 (N2875, N2860, N2138, N1740);
not NOT1 (N2876, N2844);
not NOT1 (N2877, N2865);
buf BUF1 (N2878, N2849);
not NOT1 (N2879, N2878);
nor NOR4 (N2880, N2873, N1479, N2565, N1129);
and AND2 (N2881, N2867, N1676);
and AND3 (N2882, N2846, N1982, N1484);
or OR4 (N2883, N2877, N416, N231, N2319);
buf BUF1 (N2884, N2871);
nand NAND3 (N2885, N2874, N1656, N2511);
not NOT1 (N2886, N2881);
nor NOR3 (N2887, N2885, N865, N52);
xor XOR2 (N2888, N2884, N1679);
nand NAND3 (N2889, N2882, N1544, N2459);
or OR4 (N2890, N2886, N1676, N1717, N151);
not NOT1 (N2891, N2880);
nand NAND4 (N2892, N2889, N2165, N58, N1392);
not NOT1 (N2893, N2891);
nor NOR3 (N2894, N2892, N2845, N2310);
buf BUF1 (N2895, N2888);
nor NOR4 (N2896, N2890, N97, N598, N1319);
and AND2 (N2897, N2887, N1678);
not NOT1 (N2898, N2883);
and AND3 (N2899, N2872, N665, N2818);
xor XOR2 (N2900, N2893, N1895);
not NOT1 (N2901, N2898);
buf BUF1 (N2902, N2876);
or OR2 (N2903, N2895, N2342);
buf BUF1 (N2904, N2899);
xor XOR2 (N2905, N2894, N100);
and AND3 (N2906, N2902, N1475, N2628);
buf BUF1 (N2907, N2875);
nand NAND3 (N2908, N2907, N1257, N2012);
nor NOR4 (N2909, N2908, N953, N1025, N492);
buf BUF1 (N2910, N2897);
or OR2 (N2911, N2905, N1187);
or OR2 (N2912, N2900, N1573);
not NOT1 (N2913, N2910);
nor NOR2 (N2914, N2913, N2540);
and AND4 (N2915, N2896, N1913, N2367, N2792);
not NOT1 (N2916, N2879);
nand NAND3 (N2917, N2914, N2347, N1463);
xor XOR2 (N2918, N2916, N969);
and AND3 (N2919, N2901, N1478, N1675);
buf BUF1 (N2920, N2909);
and AND2 (N2921, N2919, N790);
or OR4 (N2922, N2912, N205, N2393, N1526);
nor NOR2 (N2923, N2903, N2528);
and AND2 (N2924, N2906, N2859);
or OR2 (N2925, N2922, N1710);
and AND4 (N2926, N2904, N335, N2169, N861);
xor XOR2 (N2927, N2917, N407);
xor XOR2 (N2928, N2920, N2650);
not NOT1 (N2929, N2927);
xor XOR2 (N2930, N2928, N1907);
not NOT1 (N2931, N2926);
xor XOR2 (N2932, N2915, N2308);
not NOT1 (N2933, N2921);
or OR2 (N2934, N2930, N2614);
buf BUF1 (N2935, N2911);
buf BUF1 (N2936, N2931);
buf BUF1 (N2937, N2925);
nor NOR2 (N2938, N2933, N2730);
or OR4 (N2939, N2938, N1604, N1412, N2101);
not NOT1 (N2940, N2937);
nand NAND3 (N2941, N2934, N1114, N1603);
or OR3 (N2942, N2918, N2687, N2293);
and AND4 (N2943, N2942, N1185, N2911, N2228);
nor NOR3 (N2944, N2939, N2440, N2307);
buf BUF1 (N2945, N2940);
nor NOR2 (N2946, N2924, N2889);
or OR2 (N2947, N2944, N2799);
xor XOR2 (N2948, N2947, N2269);
nor NOR3 (N2949, N2946, N1525, N2928);
nand NAND3 (N2950, N2936, N2187, N2240);
buf BUF1 (N2951, N2943);
nor NOR3 (N2952, N2950, N1384, N960);
nor NOR4 (N2953, N2923, N27, N2538, N601);
and AND2 (N2954, N2951, N2421);
or OR2 (N2955, N2932, N2851);
or OR4 (N2956, N2954, N1175, N1941, N1427);
buf BUF1 (N2957, N2955);
not NOT1 (N2958, N2953);
and AND2 (N2959, N2929, N2494);
buf BUF1 (N2960, N2949);
nand NAND3 (N2961, N2957, N310, N32);
xor XOR2 (N2962, N2961, N2783);
nor NOR2 (N2963, N2962, N2575);
not NOT1 (N2964, N2952);
buf BUF1 (N2965, N2964);
nand NAND3 (N2966, N2965, N2591, N46);
nand NAND2 (N2967, N2966, N1081);
or OR2 (N2968, N2945, N1306);
or OR3 (N2969, N2948, N1481, N2210);
nor NOR4 (N2970, N2956, N1540, N2203, N1465);
xor XOR2 (N2971, N2970, N2548);
xor XOR2 (N2972, N2967, N2009);
buf BUF1 (N2973, N2971);
not NOT1 (N2974, N2941);
nor NOR2 (N2975, N2963, N1246);
and AND3 (N2976, N2935, N2565, N1138);
and AND2 (N2977, N2972, N2414);
xor XOR2 (N2978, N2975, N2211);
xor XOR2 (N2979, N2974, N87);
and AND3 (N2980, N2969, N78, N1148);
not NOT1 (N2981, N2976);
nand NAND2 (N2982, N2981, N2973);
and AND2 (N2983, N374, N1091);
or OR2 (N2984, N2979, N1353);
or OR4 (N2985, N2977, N2064, N2590, N982);
or OR3 (N2986, N2984, N2652, N2832);
or OR2 (N2987, N2959, N920);
nor NOR4 (N2988, N2980, N554, N611, N1952);
nor NOR4 (N2989, N2985, N834, N1549, N2345);
nand NAND3 (N2990, N2989, N2319, N854);
not NOT1 (N2991, N2986);
nand NAND4 (N2992, N2968, N1473, N2648, N1458);
nand NAND4 (N2993, N2988, N551, N1829, N121);
nor NOR4 (N2994, N2992, N800, N413, N61);
buf BUF1 (N2995, N2960);
nand NAND2 (N2996, N2958, N2937);
xor XOR2 (N2997, N2982, N468);
or OR2 (N2998, N2997, N847);
xor XOR2 (N2999, N2998, N1393);
and AND2 (N3000, N2987, N1577);
not NOT1 (N3001, N2983);
and AND4 (N3002, N2999, N1359, N1625, N1685);
or OR3 (N3003, N3001, N1378, N200);
xor XOR2 (N3004, N2991, N856);
not NOT1 (N3005, N2978);
nor NOR4 (N3006, N2995, N1678, N428, N95);
nand NAND4 (N3007, N3000, N2617, N2668, N1224);
nor NOR2 (N3008, N2990, N548);
or OR2 (N3009, N3005, N602);
and AND4 (N3010, N2994, N555, N2854, N314);
nor NOR2 (N3011, N3007, N1488);
and AND3 (N3012, N3006, N348, N734);
and AND3 (N3013, N3008, N2244, N1766);
or OR2 (N3014, N2996, N2937);
xor XOR2 (N3015, N3010, N2100);
not NOT1 (N3016, N3002);
nor NOR3 (N3017, N3004, N1441, N1023);
and AND4 (N3018, N3009, N2273, N1072, N2808);
buf BUF1 (N3019, N3016);
nand NAND2 (N3020, N3014, N2771);
buf BUF1 (N3021, N3020);
nor NOR4 (N3022, N2993, N793, N1710, N807);
or OR3 (N3023, N3022, N2811, N1565);
and AND2 (N3024, N3018, N1634);
and AND3 (N3025, N3015, N3002, N518);
not NOT1 (N3026, N3021);
or OR3 (N3027, N3024, N2181, N2205);
xor XOR2 (N3028, N3026, N2767);
xor XOR2 (N3029, N3003, N1183);
and AND4 (N3030, N3025, N946, N2201, N2252);
nor NOR3 (N3031, N3017, N2677, N710);
or OR4 (N3032, N3023, N172, N2634, N2456);
or OR3 (N3033, N3031, N1323, N1989);
buf BUF1 (N3034, N3033);
buf BUF1 (N3035, N3013);
xor XOR2 (N3036, N3029, N2281);
and AND4 (N3037, N3027, N2055, N733, N1376);
and AND3 (N3038, N3028, N1794, N2551);
buf BUF1 (N3039, N3011);
and AND2 (N3040, N3032, N1895);
and AND4 (N3041, N3019, N2419, N319, N547);
not NOT1 (N3042, N3038);
and AND2 (N3043, N3036, N267);
nor NOR2 (N3044, N3040, N864);
xor XOR2 (N3045, N3035, N1435);
nor NOR3 (N3046, N3012, N164, N21);
nand NAND2 (N3047, N3037, N1817);
not NOT1 (N3048, N3044);
and AND3 (N3049, N3039, N1680, N1601);
not NOT1 (N3050, N3034);
or OR2 (N3051, N3047, N656);
xor XOR2 (N3052, N3041, N2894);
buf BUF1 (N3053, N3046);
and AND2 (N3054, N3045, N2190);
nand NAND2 (N3055, N3043, N727);
not NOT1 (N3056, N3030);
nand NAND4 (N3057, N3054, N1087, N1994, N1387);
buf BUF1 (N3058, N3049);
xor XOR2 (N3059, N3042, N1624);
xor XOR2 (N3060, N3048, N2591);
or OR4 (N3061, N3060, N284, N2688, N2627);
not NOT1 (N3062, N3056);
or OR2 (N3063, N3058, N1845);
not NOT1 (N3064, N3061);
xor XOR2 (N3065, N3050, N2376);
nand NAND2 (N3066, N3063, N1270);
not NOT1 (N3067, N3055);
buf BUF1 (N3068, N3052);
xor XOR2 (N3069, N3064, N1290);
and AND2 (N3070, N3057, N2993);
buf BUF1 (N3071, N3059);
or OR3 (N3072, N3070, N2513, N2283);
nand NAND4 (N3073, N3065, N1957, N356, N1100);
nor NOR2 (N3074, N3071, N3037);
nand NAND4 (N3075, N3051, N517, N1223, N2730);
nand NAND2 (N3076, N3068, N2935);
or OR4 (N3077, N3053, N245, N1444, N1488);
buf BUF1 (N3078, N3069);
not NOT1 (N3079, N3066);
nor NOR4 (N3080, N3079, N2169, N2648, N213);
xor XOR2 (N3081, N3073, N2196);
buf BUF1 (N3082, N3075);
not NOT1 (N3083, N3074);
nor NOR2 (N3084, N3067, N1930);
nor NOR4 (N3085, N3080, N27, N1558, N1029);
xor XOR2 (N3086, N3078, N1004);
xor XOR2 (N3087, N3083, N1985);
or OR3 (N3088, N3072, N2292, N3061);
or OR3 (N3089, N3087, N1778, N2013);
xor XOR2 (N3090, N3082, N1691);
not NOT1 (N3091, N3088);
or OR4 (N3092, N3084, N1917, N270, N1357);
nor NOR3 (N3093, N3090, N467, N2274);
buf BUF1 (N3094, N3081);
xor XOR2 (N3095, N3077, N2454);
and AND3 (N3096, N3089, N480, N160);
nand NAND2 (N3097, N3091, N2623);
nor NOR3 (N3098, N3092, N1247, N1890);
or OR2 (N3099, N3094, N628);
xor XOR2 (N3100, N3076, N2821);
nor NOR4 (N3101, N3098, N1276, N2332, N2446);
or OR3 (N3102, N3093, N40, N886);
and AND3 (N3103, N3096, N1311, N2698);
or OR3 (N3104, N3062, N1994, N2754);
nand NAND4 (N3105, N3102, N831, N1319, N2967);
nand NAND2 (N3106, N3103, N1409);
nand NAND2 (N3107, N3100, N256);
buf BUF1 (N3108, N3085);
nand NAND2 (N3109, N3095, N2130);
buf BUF1 (N3110, N3106);
nor NOR3 (N3111, N3101, N1360, N2831);
xor XOR2 (N3112, N3107, N1316);
nand NAND2 (N3113, N3097, N3095);
nor NOR2 (N3114, N3112, N2283);
or OR3 (N3115, N3108, N2976, N2159);
nor NOR2 (N3116, N3099, N131);
and AND3 (N3117, N3105, N1984, N2482);
xor XOR2 (N3118, N3109, N2892);
buf BUF1 (N3119, N3114);
nand NAND3 (N3120, N3119, N2825, N2725);
or OR3 (N3121, N3120, N639, N2674);
buf BUF1 (N3122, N3115);
and AND4 (N3123, N3118, N1736, N2787, N2549);
or OR2 (N3124, N3113, N1259);
xor XOR2 (N3125, N3117, N870);
or OR2 (N3126, N3123, N2498);
buf BUF1 (N3127, N3116);
and AND2 (N3128, N3086, N1665);
nand NAND2 (N3129, N3110, N2175);
or OR2 (N3130, N3122, N22);
nor NOR2 (N3131, N3126, N873);
buf BUF1 (N3132, N3129);
buf BUF1 (N3133, N3121);
buf BUF1 (N3134, N3131);
or OR3 (N3135, N3132, N2143, N2294);
xor XOR2 (N3136, N3128, N592);
and AND3 (N3137, N3135, N1571, N2704);
not NOT1 (N3138, N3127);
and AND2 (N3139, N3137, N1866);
and AND4 (N3140, N3111, N45, N2922, N645);
nand NAND3 (N3141, N3138, N834, N2633);
nand NAND3 (N3142, N3130, N2670, N2026);
not NOT1 (N3143, N3139);
nand NAND2 (N3144, N3125, N2803);
and AND2 (N3145, N3134, N1369);
xor XOR2 (N3146, N3104, N60);
xor XOR2 (N3147, N3140, N2362);
and AND3 (N3148, N3142, N2233, N1206);
and AND3 (N3149, N3143, N513, N1530);
nor NOR2 (N3150, N3148, N453);
xor XOR2 (N3151, N3144, N982);
nand NAND4 (N3152, N3147, N2362, N2116, N2911);
not NOT1 (N3153, N3152);
not NOT1 (N3154, N3153);
not NOT1 (N3155, N3146);
nand NAND3 (N3156, N3151, N3024, N973);
or OR2 (N3157, N3154, N204);
or OR3 (N3158, N3133, N267, N2264);
nand NAND2 (N3159, N3136, N1212);
nand NAND3 (N3160, N3158, N2299, N125);
buf BUF1 (N3161, N3149);
xor XOR2 (N3162, N3161, N1805);
xor XOR2 (N3163, N3160, N554);
and AND4 (N3164, N3150, N2840, N2154, N270);
nand NAND2 (N3165, N3145, N1376);
and AND4 (N3166, N3141, N2205, N2485, N2105);
not NOT1 (N3167, N3155);
not NOT1 (N3168, N3159);
not NOT1 (N3169, N3156);
and AND4 (N3170, N3165, N1135, N732, N1951);
or OR2 (N3171, N3170, N302);
nand NAND4 (N3172, N3168, N2416, N2313, N1251);
not NOT1 (N3173, N3167);
and AND2 (N3174, N3164, N2913);
not NOT1 (N3175, N3169);
not NOT1 (N3176, N3171);
not NOT1 (N3177, N3163);
buf BUF1 (N3178, N3172);
not NOT1 (N3179, N3175);
and AND3 (N3180, N3174, N2352, N2724);
or OR3 (N3181, N3124, N1981, N3176);
or OR4 (N3182, N1612, N1411, N1660, N2905);
and AND4 (N3183, N3162, N854, N2950, N3056);
or OR4 (N3184, N3178, N113, N236, N3026);
and AND2 (N3185, N3157, N1138);
not NOT1 (N3186, N3183);
or OR3 (N3187, N3185, N2294, N2830);
xor XOR2 (N3188, N3180, N1286);
or OR2 (N3189, N3187, N2708);
and AND2 (N3190, N3182, N396);
not NOT1 (N3191, N3190);
or OR4 (N3192, N3166, N2812, N2266, N91);
and AND4 (N3193, N3173, N1516, N2424, N2996);
or OR3 (N3194, N3193, N1269, N1055);
not NOT1 (N3195, N3181);
nor NOR2 (N3196, N3189, N3147);
or OR4 (N3197, N3192, N2525, N575, N2343);
nand NAND3 (N3198, N3186, N1459, N2720);
nor NOR3 (N3199, N3177, N2334, N1475);
or OR3 (N3200, N3196, N3188, N656);
or OR2 (N3201, N2432, N2873);
not NOT1 (N3202, N3200);
xor XOR2 (N3203, N3202, N585);
nor NOR4 (N3204, N3198, N1718, N487, N1467);
nor NOR4 (N3205, N3191, N1206, N54, N3191);
buf BUF1 (N3206, N3194);
not NOT1 (N3207, N3203);
not NOT1 (N3208, N3205);
nor NOR3 (N3209, N3204, N686, N1142);
or OR4 (N3210, N3195, N913, N2997, N2339);
buf BUF1 (N3211, N3199);
nand NAND3 (N3212, N3208, N1432, N1079);
nor NOR3 (N3213, N3179, N3018, N2214);
xor XOR2 (N3214, N3207, N1353);
or OR4 (N3215, N3209, N2972, N509, N2636);
xor XOR2 (N3216, N3213, N3051);
nor NOR4 (N3217, N3215, N131, N901, N2917);
not NOT1 (N3218, N3217);
not NOT1 (N3219, N3216);
xor XOR2 (N3220, N3210, N2475);
or OR4 (N3221, N3214, N259, N2044, N1014);
nand NAND4 (N3222, N3211, N1476, N1043, N291);
nand NAND3 (N3223, N3197, N523, N1406);
not NOT1 (N3224, N3218);
xor XOR2 (N3225, N3224, N1404);
not NOT1 (N3226, N3184);
xor XOR2 (N3227, N3222, N1259);
xor XOR2 (N3228, N3220, N1150);
not NOT1 (N3229, N3227);
or OR4 (N3230, N3226, N2213, N746, N2748);
not NOT1 (N3231, N3219);
or OR2 (N3232, N3206, N2570);
or OR3 (N3233, N3212, N2698, N2169);
nor NOR3 (N3234, N3223, N3131, N1151);
and AND4 (N3235, N3230, N2402, N2939, N1579);
or OR2 (N3236, N3225, N985);
nor NOR3 (N3237, N3229, N190, N215);
xor XOR2 (N3238, N3233, N1594);
not NOT1 (N3239, N3235);
nand NAND2 (N3240, N3237, N376);
not NOT1 (N3241, N3228);
buf BUF1 (N3242, N3232);
xor XOR2 (N3243, N3242, N1750);
nand NAND2 (N3244, N3239, N3099);
nand NAND3 (N3245, N3201, N2436, N88);
not NOT1 (N3246, N3238);
or OR2 (N3247, N3244, N1188);
xor XOR2 (N3248, N3243, N1594);
and AND3 (N3249, N3236, N1898, N3240);
nor NOR3 (N3250, N1707, N3099, N3050);
xor XOR2 (N3251, N3231, N316);
buf BUF1 (N3252, N3234);
nor NOR3 (N3253, N3241, N1688, N3052);
nand NAND3 (N3254, N3247, N2091, N1027);
nand NAND2 (N3255, N3246, N2601);
and AND4 (N3256, N3254, N1475, N2208, N2843);
buf BUF1 (N3257, N3249);
and AND3 (N3258, N3256, N2120, N473);
buf BUF1 (N3259, N3250);
nand NAND2 (N3260, N3258, N1161);
not NOT1 (N3261, N3221);
and AND4 (N3262, N3251, N2393, N1595, N1511);
not NOT1 (N3263, N3253);
or OR3 (N3264, N3255, N2592, N1926);
nor NOR4 (N3265, N3263, N2491, N2236, N3132);
and AND2 (N3266, N3248, N417);
not NOT1 (N3267, N3262);
not NOT1 (N3268, N3264);
or OR2 (N3269, N3245, N2050);
or OR4 (N3270, N3268, N195, N370, N996);
and AND4 (N3271, N3261, N2368, N1294, N1396);
nand NAND4 (N3272, N3265, N2391, N2458, N118);
or OR4 (N3273, N3260, N2074, N1011, N2087);
nor NOR2 (N3274, N3267, N167);
nand NAND2 (N3275, N3273, N94);
not NOT1 (N3276, N3266);
and AND3 (N3277, N3275, N3174, N359);
nor NOR3 (N3278, N3257, N1660, N1320);
not NOT1 (N3279, N3252);
not NOT1 (N3280, N3272);
xor XOR2 (N3281, N3279, N646);
not NOT1 (N3282, N3276);
buf BUF1 (N3283, N3270);
buf BUF1 (N3284, N3259);
not NOT1 (N3285, N3284);
and AND4 (N3286, N3278, N897, N2745, N2889);
not NOT1 (N3287, N3269);
and AND2 (N3288, N3282, N1371);
nand NAND2 (N3289, N3274, N693);
or OR4 (N3290, N3288, N2383, N1034, N2776);
or OR4 (N3291, N3290, N1260, N2411, N1436);
nor NOR4 (N3292, N3287, N1944, N2546, N2188);
xor XOR2 (N3293, N3280, N2372);
or OR2 (N3294, N3293, N315);
or OR4 (N3295, N3277, N705, N3208, N2150);
nand NAND3 (N3296, N3285, N2604, N846);
nand NAND2 (N3297, N3296, N3039);
buf BUF1 (N3298, N3291);
nor NOR4 (N3299, N3286, N1252, N3194, N1682);
nor NOR2 (N3300, N3294, N1784);
buf BUF1 (N3301, N3299);
xor XOR2 (N3302, N3283, N300);
nor NOR4 (N3303, N3298, N2672, N3192, N1844);
nor NOR3 (N3304, N3271, N2311, N804);
or OR3 (N3305, N3300, N654, N1218);
buf BUF1 (N3306, N3295);
xor XOR2 (N3307, N3306, N1526);
nor NOR3 (N3308, N3303, N845, N3227);
nand NAND2 (N3309, N3281, N1958);
nor NOR4 (N3310, N3305, N2332, N2936, N1603);
buf BUF1 (N3311, N3304);
not NOT1 (N3312, N3292);
nand NAND3 (N3313, N3289, N253, N1153);
not NOT1 (N3314, N3307);
and AND4 (N3315, N3297, N2515, N1798, N1605);
and AND4 (N3316, N3309, N2054, N1646, N1901);
not NOT1 (N3317, N3314);
or OR3 (N3318, N3308, N1463, N1505);
not NOT1 (N3319, N3315);
buf BUF1 (N3320, N3301);
or OR4 (N3321, N3312, N269, N571, N94);
not NOT1 (N3322, N3317);
nor NOR4 (N3323, N3311, N860, N330, N1061);
nor NOR3 (N3324, N3313, N444, N1648);
or OR4 (N3325, N3310, N527, N1416, N553);
xor XOR2 (N3326, N3320, N2251);
xor XOR2 (N3327, N3323, N61);
nor NOR3 (N3328, N3316, N2340, N3247);
not NOT1 (N3329, N3321);
xor XOR2 (N3330, N3302, N450);
buf BUF1 (N3331, N3327);
not NOT1 (N3332, N3322);
buf BUF1 (N3333, N3325);
nand NAND4 (N3334, N3331, N1434, N34, N1900);
nand NAND2 (N3335, N3333, N1195);
not NOT1 (N3336, N3324);
and AND3 (N3337, N3319, N1094, N1176);
not NOT1 (N3338, N3336);
buf BUF1 (N3339, N3332);
nor NOR4 (N3340, N3326, N337, N2726, N2048);
and AND2 (N3341, N3339, N2532);
xor XOR2 (N3342, N3334, N2016);
or OR3 (N3343, N3329, N272, N1859);
nor NOR2 (N3344, N3318, N1356);
buf BUF1 (N3345, N3341);
xor XOR2 (N3346, N3328, N2775);
and AND3 (N3347, N3340, N1002, N2193);
xor XOR2 (N3348, N3342, N1775);
not NOT1 (N3349, N3347);
nor NOR2 (N3350, N3349, N2572);
xor XOR2 (N3351, N3330, N2636);
and AND3 (N3352, N3343, N3007, N2582);
buf BUF1 (N3353, N3346);
not NOT1 (N3354, N3352);
nand NAND2 (N3355, N3335, N2894);
buf BUF1 (N3356, N3344);
nor NOR4 (N3357, N3353, N2881, N2136, N1329);
and AND3 (N3358, N3348, N606, N991);
xor XOR2 (N3359, N3337, N282);
buf BUF1 (N3360, N3357);
and AND3 (N3361, N3358, N3157, N3086);
not NOT1 (N3362, N3361);
buf BUF1 (N3363, N3345);
buf BUF1 (N3364, N3362);
xor XOR2 (N3365, N3363, N2830);
buf BUF1 (N3366, N3350);
or OR3 (N3367, N3364, N378, N2320);
nor NOR3 (N3368, N3366, N624, N2060);
and AND4 (N3369, N3356, N2014, N1726, N2234);
xor XOR2 (N3370, N3359, N338);
nor NOR2 (N3371, N3355, N2111);
nor NOR4 (N3372, N3354, N128, N408, N61);
or OR3 (N3373, N3360, N160, N2388);
or OR2 (N3374, N3369, N859);
buf BUF1 (N3375, N3351);
nand NAND4 (N3376, N3370, N490, N1007, N1138);
not NOT1 (N3377, N3374);
and AND2 (N3378, N3365, N573);
or OR4 (N3379, N3368, N2437, N1231, N2202);
nor NOR3 (N3380, N3367, N645, N2873);
and AND4 (N3381, N3371, N1267, N451, N1788);
buf BUF1 (N3382, N3381);
not NOT1 (N3383, N3379);
and AND4 (N3384, N3373, N2947, N1074, N436);
not NOT1 (N3385, N3377);
not NOT1 (N3386, N3376);
xor XOR2 (N3387, N3384, N2241);
or OR4 (N3388, N3372, N2216, N3112, N180);
and AND2 (N3389, N3385, N2266);
not NOT1 (N3390, N3378);
and AND2 (N3391, N3390, N2201);
nor NOR4 (N3392, N3389, N42, N3151, N3380);
buf BUF1 (N3393, N2438);
nor NOR3 (N3394, N3382, N2207, N2152);
xor XOR2 (N3395, N3387, N2321);
and AND3 (N3396, N3386, N3351, N2610);
nand NAND4 (N3397, N3375, N1941, N2604, N2885);
nand NAND3 (N3398, N3396, N378, N904);
or OR3 (N3399, N3392, N2322, N1280);
nand NAND3 (N3400, N3393, N3036, N1449);
xor XOR2 (N3401, N3388, N2508);
buf BUF1 (N3402, N3400);
not NOT1 (N3403, N3402);
or OR3 (N3404, N3403, N1752, N2090);
xor XOR2 (N3405, N3397, N126);
xor XOR2 (N3406, N3391, N1130);
xor XOR2 (N3407, N3395, N1549);
or OR2 (N3408, N3398, N1082);
nand NAND2 (N3409, N3394, N2399);
and AND4 (N3410, N3407, N1856, N2884, N924);
nor NOR2 (N3411, N3405, N1686);
nand NAND3 (N3412, N3383, N2437, N929);
nor NOR4 (N3413, N3404, N596, N2058, N253);
nor NOR2 (N3414, N3409, N752);
not NOT1 (N3415, N3413);
and AND4 (N3416, N3414, N2314, N1112, N1434);
or OR2 (N3417, N3410, N3174);
and AND2 (N3418, N3406, N2259);
and AND4 (N3419, N3401, N2435, N3046, N1543);
nand NAND2 (N3420, N3419, N2461);
xor XOR2 (N3421, N3420, N417);
or OR2 (N3422, N3417, N1044);
buf BUF1 (N3423, N3422);
buf BUF1 (N3424, N3421);
not NOT1 (N3425, N3416);
xor XOR2 (N3426, N3408, N338);
nor NOR3 (N3427, N3399, N883, N2161);
and AND2 (N3428, N3423, N219);
xor XOR2 (N3429, N3418, N1045);
and AND3 (N3430, N3428, N2968, N637);
or OR3 (N3431, N3425, N1395, N1165);
not NOT1 (N3432, N3415);
and AND3 (N3433, N3427, N829, N2468);
not NOT1 (N3434, N3426);
nand NAND2 (N3435, N3412, N2131);
or OR4 (N3436, N3429, N697, N3407, N1650);
buf BUF1 (N3437, N3338);
or OR4 (N3438, N3436, N2524, N1872, N2759);
nand NAND3 (N3439, N3424, N2894, N859);
buf BUF1 (N3440, N3435);
nand NAND2 (N3441, N3440, N2022);
xor XOR2 (N3442, N3438, N1706);
not NOT1 (N3443, N3430);
buf BUF1 (N3444, N3443);
nand NAND3 (N3445, N3441, N2778, N1050);
nand NAND4 (N3446, N3439, N1176, N503, N3438);
not NOT1 (N3447, N3411);
xor XOR2 (N3448, N3437, N2906);
and AND4 (N3449, N3446, N2064, N1575, N1166);
or OR2 (N3450, N3447, N1949);
nand NAND4 (N3451, N3450, N1213, N3002, N2288);
nor NOR4 (N3452, N3431, N2773, N1845, N473);
or OR2 (N3453, N3444, N252);
nor NOR4 (N3454, N3453, N134, N2589, N2198);
not NOT1 (N3455, N3442);
nor NOR4 (N3456, N3434, N2234, N2050, N1891);
not NOT1 (N3457, N3445);
nor NOR3 (N3458, N3448, N902, N2410);
or OR2 (N3459, N3449, N1503);
not NOT1 (N3460, N3454);
nand NAND4 (N3461, N3452, N3181, N1457, N2042);
buf BUF1 (N3462, N3459);
or OR3 (N3463, N3455, N1598, N440);
xor XOR2 (N3464, N3461, N32);
nand NAND3 (N3465, N3432, N1568, N93);
xor XOR2 (N3466, N3457, N1589);
nor NOR2 (N3467, N3451, N876);
nand NAND2 (N3468, N3464, N1142);
and AND2 (N3469, N3468, N1681);
buf BUF1 (N3470, N3465);
nor NOR4 (N3471, N3460, N3034, N3167, N1393);
or OR4 (N3472, N3470, N2144, N1406, N2237);
nor NOR2 (N3473, N3467, N566);
nand NAND2 (N3474, N3471, N224);
xor XOR2 (N3475, N3458, N1762);
nor NOR4 (N3476, N3433, N1233, N1996, N1127);
not NOT1 (N3477, N3474);
xor XOR2 (N3478, N3472, N1003);
buf BUF1 (N3479, N3469);
not NOT1 (N3480, N3476);
nor NOR4 (N3481, N3473, N1669, N66, N1394);
and AND3 (N3482, N3477, N2667, N3478);
and AND3 (N3483, N3216, N867, N1649);
xor XOR2 (N3484, N3466, N747);
buf BUF1 (N3485, N3462);
not NOT1 (N3486, N3481);
or OR4 (N3487, N3475, N1712, N2406, N1456);
nor NOR2 (N3488, N3463, N3210);
and AND3 (N3489, N3486, N314, N1626);
and AND2 (N3490, N3483, N1905);
nand NAND2 (N3491, N3487, N1797);
buf BUF1 (N3492, N3484);
not NOT1 (N3493, N3482);
buf BUF1 (N3494, N3492);
nor NOR3 (N3495, N3456, N3153, N563);
or OR4 (N3496, N3479, N2318, N1031, N2875);
xor XOR2 (N3497, N3485, N1669);
not NOT1 (N3498, N3497);
xor XOR2 (N3499, N3496, N1863);
not NOT1 (N3500, N3480);
buf BUF1 (N3501, N3491);
not NOT1 (N3502, N3490);
nor NOR2 (N3503, N3500, N3379);
and AND3 (N3504, N3501, N1636, N3375);
xor XOR2 (N3505, N3503, N1150);
xor XOR2 (N3506, N3505, N2002);
buf BUF1 (N3507, N3495);
or OR2 (N3508, N3493, N2772);
nor NOR3 (N3509, N3506, N2079, N178);
not NOT1 (N3510, N3504);
or OR3 (N3511, N3508, N1903, N1033);
not NOT1 (N3512, N3507);
buf BUF1 (N3513, N3489);
or OR2 (N3514, N3512, N1910);
or OR3 (N3515, N3513, N924, N1508);
nor NOR4 (N3516, N3510, N1704, N257, N615);
and AND2 (N3517, N3516, N1337);
and AND2 (N3518, N3514, N1943);
buf BUF1 (N3519, N3511);
or OR3 (N3520, N3502, N3420, N1046);
and AND2 (N3521, N3515, N2935);
or OR3 (N3522, N3509, N156, N1258);
nand NAND3 (N3523, N3520, N3443, N3058);
xor XOR2 (N3524, N3519, N702);
nor NOR3 (N3525, N3517, N2208, N3204);
or OR4 (N3526, N3498, N2851, N593, N210);
not NOT1 (N3527, N3526);
nor NOR3 (N3528, N3518, N2089, N3320);
buf BUF1 (N3529, N3525);
nand NAND3 (N3530, N3521, N2158, N1724);
nor NOR3 (N3531, N3530, N3072, N1578);
and AND4 (N3532, N3524, N3457, N2807, N2872);
nor NOR3 (N3533, N3528, N2993, N741);
nor NOR2 (N3534, N3522, N2280);
or OR3 (N3535, N3499, N632, N1526);
not NOT1 (N3536, N3532);
and AND3 (N3537, N3536, N2355, N1436);
buf BUF1 (N3538, N3535);
buf BUF1 (N3539, N3534);
or OR4 (N3540, N3527, N3438, N2514, N1963);
nor NOR3 (N3541, N3523, N154, N56);
nand NAND3 (N3542, N3541, N375, N115);
not NOT1 (N3543, N3494);
not NOT1 (N3544, N3537);
xor XOR2 (N3545, N3533, N2144);
or OR4 (N3546, N3531, N1295, N187, N2511);
xor XOR2 (N3547, N3542, N2753);
not NOT1 (N3548, N3547);
and AND3 (N3549, N3529, N2785, N164);
xor XOR2 (N3550, N3539, N2094);
or OR4 (N3551, N3488, N1085, N2139, N3335);
xor XOR2 (N3552, N3550, N3092);
or OR3 (N3553, N3544, N937, N2085);
xor XOR2 (N3554, N3546, N1738);
or OR2 (N3555, N3548, N2959);
or OR3 (N3556, N3555, N2451, N34);
xor XOR2 (N3557, N3545, N482);
buf BUF1 (N3558, N3557);
nand NAND4 (N3559, N3552, N1350, N857, N2741);
or OR2 (N3560, N3543, N2782);
nor NOR2 (N3561, N3560, N974);
xor XOR2 (N3562, N3558, N508);
nor NOR4 (N3563, N3562, N2328, N1253, N778);
and AND2 (N3564, N3559, N2595);
buf BUF1 (N3565, N3551);
and AND3 (N3566, N3563, N2873, N809);
or OR3 (N3567, N3561, N672, N2891);
not NOT1 (N3568, N3565);
or OR3 (N3569, N3556, N775, N2472);
or OR4 (N3570, N3567, N2308, N1223, N596);
nor NOR3 (N3571, N3538, N1278, N769);
nor NOR2 (N3572, N3568, N2287);
and AND3 (N3573, N3572, N872, N1579);
nor NOR3 (N3574, N3570, N1674, N1620);
buf BUF1 (N3575, N3573);
nand NAND3 (N3576, N3571, N432, N276);
and AND2 (N3577, N3566, N1289);
not NOT1 (N3578, N3554);
nand NAND2 (N3579, N3577, N1255);
xor XOR2 (N3580, N3575, N2245);
nor NOR2 (N3581, N3549, N1369);
nor NOR4 (N3582, N3578, N917, N2345, N1666);
xor XOR2 (N3583, N3574, N963);
nor NOR3 (N3584, N3580, N1200, N2287);
buf BUF1 (N3585, N3583);
nor NOR3 (N3586, N3582, N2739, N3090);
buf BUF1 (N3587, N3586);
or OR4 (N3588, N3579, N1363, N3315, N3155);
buf BUF1 (N3589, N3588);
nor NOR2 (N3590, N3540, N2491);
and AND2 (N3591, N3569, N1642);
nand NAND3 (N3592, N3581, N987, N3050);
or OR3 (N3593, N3587, N2779, N998);
and AND2 (N3594, N3593, N3517);
nand NAND2 (N3595, N3585, N2883);
xor XOR2 (N3596, N3592, N3028);
xor XOR2 (N3597, N3564, N3178);
nand NAND4 (N3598, N3584, N86, N468, N3278);
not NOT1 (N3599, N3597);
xor XOR2 (N3600, N3594, N189);
xor XOR2 (N3601, N3576, N1487);
xor XOR2 (N3602, N3599, N236);
nor NOR2 (N3603, N3590, N1859);
nor NOR2 (N3604, N3602, N1016);
nand NAND3 (N3605, N3589, N109, N943);
buf BUF1 (N3606, N3591);
xor XOR2 (N3607, N3596, N158);
nand NAND3 (N3608, N3601, N183, N275);
nor NOR4 (N3609, N3598, N1859, N801, N2063);
buf BUF1 (N3610, N3606);
not NOT1 (N3611, N3603);
nor NOR4 (N3612, N3605, N3456, N21, N1709);
xor XOR2 (N3613, N3610, N2027);
buf BUF1 (N3614, N3595);
nor NOR2 (N3615, N3613, N1611);
nor NOR2 (N3616, N3615, N1018);
buf BUF1 (N3617, N3608);
buf BUF1 (N3618, N3553);
xor XOR2 (N3619, N3616, N1119);
and AND3 (N3620, N3617, N2207, N55);
nor NOR4 (N3621, N3614, N3054, N3216, N737);
nand NAND2 (N3622, N3619, N1387);
buf BUF1 (N3623, N3620);
xor XOR2 (N3624, N3621, N63);
nand NAND2 (N3625, N3618, N3300);
nor NOR4 (N3626, N3622, N1816, N2931, N903);
xor XOR2 (N3627, N3625, N3063);
buf BUF1 (N3628, N3626);
not NOT1 (N3629, N3604);
xor XOR2 (N3630, N3628, N1755);
nand NAND4 (N3631, N3630, N1583, N1228, N2309);
or OR2 (N3632, N3629, N3592);
nand NAND4 (N3633, N3609, N404, N1707, N642);
not NOT1 (N3634, N3600);
not NOT1 (N3635, N3633);
buf BUF1 (N3636, N3611);
xor XOR2 (N3637, N3636, N1618);
nor NOR2 (N3638, N3635, N998);
xor XOR2 (N3639, N3631, N3355);
nor NOR2 (N3640, N3624, N676);
xor XOR2 (N3641, N3632, N384);
or OR4 (N3642, N3612, N1930, N3136, N339);
nor NOR4 (N3643, N3637, N3065, N1612, N2997);
nor NOR4 (N3644, N3638, N2508, N1941, N507);
buf BUF1 (N3645, N3634);
or OR4 (N3646, N3642, N3139, N505, N973);
or OR3 (N3647, N3643, N212, N1099);
not NOT1 (N3648, N3639);
xor XOR2 (N3649, N3623, N3230);
nor NOR2 (N3650, N3627, N3197);
not NOT1 (N3651, N3645);
or OR4 (N3652, N3647, N658, N798, N2606);
xor XOR2 (N3653, N3607, N1210);
nand NAND2 (N3654, N3653, N1442);
xor XOR2 (N3655, N3652, N137);
or OR2 (N3656, N3646, N986);
nor NOR4 (N3657, N3651, N1771, N2181, N2124);
nor NOR3 (N3658, N3654, N2087, N867);
and AND2 (N3659, N3648, N680);
not NOT1 (N3660, N3640);
and AND3 (N3661, N3658, N1278, N3452);
nand NAND2 (N3662, N3657, N1190);
nand NAND2 (N3663, N3659, N242);
and AND3 (N3664, N3641, N2449, N1686);
xor XOR2 (N3665, N3661, N3334);
nand NAND2 (N3666, N3665, N2944);
not NOT1 (N3667, N3663);
or OR3 (N3668, N3666, N536, N3191);
buf BUF1 (N3669, N3662);
or OR4 (N3670, N3649, N528, N1789, N3540);
nand NAND4 (N3671, N3644, N2847, N2436, N2411);
and AND2 (N3672, N3655, N37);
or OR2 (N3673, N3656, N2026);
or OR2 (N3674, N3650, N2063);
nand NAND4 (N3675, N3660, N3254, N854, N2013);
nor NOR4 (N3676, N3670, N3557, N1979, N1587);
buf BUF1 (N3677, N3673);
nand NAND3 (N3678, N3664, N72, N2527);
and AND4 (N3679, N3671, N1945, N2739, N2373);
not NOT1 (N3680, N3676);
xor XOR2 (N3681, N3672, N2121);
or OR3 (N3682, N3675, N1142, N2940);
xor XOR2 (N3683, N3681, N1037);
nor NOR3 (N3684, N3683, N2415, N2759);
buf BUF1 (N3685, N3678);
and AND2 (N3686, N3679, N2034);
nor NOR2 (N3687, N3668, N1081);
xor XOR2 (N3688, N3685, N380);
nand NAND3 (N3689, N3684, N2232, N2336);
xor XOR2 (N3690, N3674, N1691);
nor NOR2 (N3691, N3680, N373);
xor XOR2 (N3692, N3677, N871);
not NOT1 (N3693, N3689);
xor XOR2 (N3694, N3686, N59);
nand NAND4 (N3695, N3669, N2520, N2682, N130);
nor NOR4 (N3696, N3687, N140, N611, N1788);
or OR4 (N3697, N3694, N3549, N3617, N2088);
not NOT1 (N3698, N3692);
or OR4 (N3699, N3688, N1214, N3225, N1611);
xor XOR2 (N3700, N3690, N3671);
nor NOR4 (N3701, N3696, N1615, N2806, N2795);
and AND2 (N3702, N3699, N2321);
or OR3 (N3703, N3700, N1822, N2859);
and AND3 (N3704, N3682, N3234, N3610);
xor XOR2 (N3705, N3704, N1185);
nor NOR4 (N3706, N3705, N313, N409, N1904);
xor XOR2 (N3707, N3693, N1560);
xor XOR2 (N3708, N3691, N1520);
nor NOR2 (N3709, N3706, N3075);
xor XOR2 (N3710, N3697, N2657);
nor NOR4 (N3711, N3703, N1778, N806, N2735);
nand NAND3 (N3712, N3711, N2104, N2910);
not NOT1 (N3713, N3701);
and AND2 (N3714, N3709, N681);
and AND3 (N3715, N3667, N2607, N197);
and AND2 (N3716, N3713, N2456);
or OR4 (N3717, N3695, N459, N3527, N2677);
or OR4 (N3718, N3707, N2104, N2823, N788);
nand NAND2 (N3719, N3712, N3146);
and AND4 (N3720, N3698, N2842, N917, N1946);
nor NOR4 (N3721, N3710, N3501, N1719, N3449);
and AND2 (N3722, N3716, N3682);
not NOT1 (N3723, N3718);
nand NAND3 (N3724, N3719, N998, N353);
and AND3 (N3725, N3715, N728, N283);
and AND3 (N3726, N3725, N2198, N194);
nor NOR2 (N3727, N3726, N969);
nor NOR2 (N3728, N3717, N346);
or OR4 (N3729, N3728, N2560, N1603, N969);
nand NAND2 (N3730, N3708, N265);
or OR4 (N3731, N3720, N1926, N3247, N3127);
nor NOR3 (N3732, N3730, N3293, N3389);
and AND4 (N3733, N3721, N2959, N390, N2809);
nor NOR2 (N3734, N3722, N1382);
buf BUF1 (N3735, N3724);
or OR4 (N3736, N3734, N340, N183, N3627);
nand NAND4 (N3737, N3735, N760, N2906, N532);
nor NOR4 (N3738, N3714, N2248, N616, N39);
not NOT1 (N3739, N3738);
and AND4 (N3740, N3736, N2522, N755, N3355);
nor NOR3 (N3741, N3702, N2586, N1485);
and AND2 (N3742, N3737, N555);
buf BUF1 (N3743, N3729);
not NOT1 (N3744, N3727);
and AND3 (N3745, N3742, N8, N463);
nand NAND2 (N3746, N3739, N890);
or OR3 (N3747, N3723, N718, N1446);
not NOT1 (N3748, N3731);
xor XOR2 (N3749, N3744, N217);
nor NOR3 (N3750, N3743, N2816, N3567);
nor NOR3 (N3751, N3741, N2804, N1645);
xor XOR2 (N3752, N3749, N2485);
or OR3 (N3753, N3748, N2939, N2875);
or OR4 (N3754, N3740, N613, N1215, N187);
xor XOR2 (N3755, N3745, N2732);
nor NOR3 (N3756, N3751, N2485, N845);
not NOT1 (N3757, N3747);
xor XOR2 (N3758, N3756, N689);
and AND2 (N3759, N3754, N760);
and AND3 (N3760, N3753, N1027, N3528);
not NOT1 (N3761, N3757);
and AND3 (N3762, N3761, N869, N3336);
xor XOR2 (N3763, N3760, N2473);
xor XOR2 (N3764, N3755, N3574);
buf BUF1 (N3765, N3752);
nand NAND2 (N3766, N3746, N841);
xor XOR2 (N3767, N3762, N1444);
not NOT1 (N3768, N3767);
xor XOR2 (N3769, N3763, N944);
buf BUF1 (N3770, N3732);
or OR3 (N3771, N3764, N1386, N2257);
nand NAND3 (N3772, N3768, N1621, N3535);
not NOT1 (N3773, N3770);
nand NAND4 (N3774, N3759, N64, N1797, N2366);
xor XOR2 (N3775, N3772, N782);
nor NOR4 (N3776, N3766, N1723, N970, N1664);
not NOT1 (N3777, N3733);
or OR2 (N3778, N3773, N2346);
and AND4 (N3779, N3776, N3203, N1937, N2122);
xor XOR2 (N3780, N3771, N3729);
xor XOR2 (N3781, N3765, N2648);
xor XOR2 (N3782, N3774, N3034);
or OR3 (N3783, N3781, N1372, N3707);
nand NAND4 (N3784, N3775, N1852, N3657, N1575);
or OR2 (N3785, N3758, N3544);
not NOT1 (N3786, N3769);
nor NOR2 (N3787, N3778, N446);
or OR4 (N3788, N3786, N880, N1999, N1902);
buf BUF1 (N3789, N3777);
and AND3 (N3790, N3784, N2783, N1306);
not NOT1 (N3791, N3790);
buf BUF1 (N3792, N3791);
nand NAND3 (N3793, N3779, N431, N1816);
xor XOR2 (N3794, N3789, N3040);
nor NOR4 (N3795, N3782, N672, N1260, N3766);
or OR3 (N3796, N3750, N3463, N1971);
nor NOR4 (N3797, N3787, N3215, N942, N1541);
xor XOR2 (N3798, N3792, N140);
not NOT1 (N3799, N3795);
nand NAND2 (N3800, N3785, N2325);
or OR2 (N3801, N3788, N1213);
or OR3 (N3802, N3780, N1677, N3363);
buf BUF1 (N3803, N3800);
nor NOR2 (N3804, N3801, N3710);
not NOT1 (N3805, N3796);
not NOT1 (N3806, N3803);
or OR4 (N3807, N3798, N3803, N2890, N738);
and AND2 (N3808, N3804, N2484);
buf BUF1 (N3809, N3793);
nand NAND3 (N3810, N3809, N1090, N1021);
xor XOR2 (N3811, N3805, N658);
buf BUF1 (N3812, N3810);
buf BUF1 (N3813, N3806);
nor NOR3 (N3814, N3797, N1566, N3521);
nor NOR4 (N3815, N3783, N336, N580, N1357);
nor NOR2 (N3816, N3802, N2002);
xor XOR2 (N3817, N3813, N782);
nand NAND3 (N3818, N3814, N2775, N360);
and AND2 (N3819, N3799, N2696);
xor XOR2 (N3820, N3819, N1254);
or OR3 (N3821, N3818, N2144, N1327);
or OR3 (N3822, N3820, N1707, N2232);
buf BUF1 (N3823, N3821);
and AND2 (N3824, N3815, N710);
xor XOR2 (N3825, N3812, N2786);
nand NAND3 (N3826, N3811, N3167, N1642);
nand NAND3 (N3827, N3826, N2027, N514);
and AND2 (N3828, N3807, N1639);
xor XOR2 (N3829, N3827, N2288);
and AND3 (N3830, N3817, N2241, N1905);
not NOT1 (N3831, N3829);
or OR4 (N3832, N3808, N628, N1468, N244);
or OR2 (N3833, N3831, N70);
nand NAND4 (N3834, N3833, N786, N818, N176);
nor NOR4 (N3835, N3823, N1085, N2850, N877);
xor XOR2 (N3836, N3816, N2236);
or OR2 (N3837, N3828, N1147);
buf BUF1 (N3838, N3834);
not NOT1 (N3839, N3837);
and AND4 (N3840, N3824, N1263, N1320, N788);
nor NOR2 (N3841, N3825, N2999);
and AND2 (N3842, N3839, N2567);
nand NAND4 (N3843, N3832, N3721, N1945, N1716);
and AND2 (N3844, N3838, N2871);
xor XOR2 (N3845, N3842, N3555);
or OR4 (N3846, N3830, N262, N3721, N1327);
or OR4 (N3847, N3835, N814, N294, N3121);
or OR4 (N3848, N3840, N3390, N3387, N107);
xor XOR2 (N3849, N3844, N2070);
nand NAND2 (N3850, N3849, N383);
not NOT1 (N3851, N3836);
nor NOR4 (N3852, N3851, N2255, N797, N488);
xor XOR2 (N3853, N3848, N1037);
xor XOR2 (N3854, N3850, N2810);
nand NAND4 (N3855, N3841, N1453, N1, N3126);
xor XOR2 (N3856, N3852, N447);
buf BUF1 (N3857, N3846);
buf BUF1 (N3858, N3843);
xor XOR2 (N3859, N3857, N22);
nand NAND2 (N3860, N3859, N641);
xor XOR2 (N3861, N3855, N1425);
nor NOR4 (N3862, N3861, N2521, N3510, N2822);
buf BUF1 (N3863, N3847);
buf BUF1 (N3864, N3862);
nor NOR2 (N3865, N3856, N1183);
nor NOR2 (N3866, N3794, N1115);
nand NAND4 (N3867, N3865, N2268, N1473, N3330);
or OR4 (N3868, N3858, N3862, N837, N3736);
and AND3 (N3869, N3863, N3273, N1669);
xor XOR2 (N3870, N3854, N2647);
nand NAND4 (N3871, N3864, N2057, N86, N515);
not NOT1 (N3872, N3871);
xor XOR2 (N3873, N3822, N2533);
nand NAND3 (N3874, N3869, N1152, N575);
and AND3 (N3875, N3872, N4, N133);
not NOT1 (N3876, N3853);
not NOT1 (N3877, N3875);
or OR2 (N3878, N3874, N2971);
buf BUF1 (N3879, N3867);
xor XOR2 (N3880, N3868, N3050);
and AND3 (N3881, N3879, N1158, N3680);
xor XOR2 (N3882, N3878, N716);
not NOT1 (N3883, N3881);
buf BUF1 (N3884, N3866);
and AND4 (N3885, N3845, N1927, N989, N1687);
nand NAND4 (N3886, N3873, N973, N753, N2959);
buf BUF1 (N3887, N3860);
not NOT1 (N3888, N3886);
nor NOR2 (N3889, N3870, N2685);
or OR3 (N3890, N3889, N2536, N582);
nor NOR2 (N3891, N3888, N743);
nand NAND4 (N3892, N3885, N3672, N817, N312);
xor XOR2 (N3893, N3884, N1693);
not NOT1 (N3894, N3890);
buf BUF1 (N3895, N3891);
or OR2 (N3896, N3882, N3328);
nand NAND2 (N3897, N3876, N447);
not NOT1 (N3898, N3896);
buf BUF1 (N3899, N3883);
nand NAND3 (N3900, N3899, N1250, N347);
nand NAND2 (N3901, N3900, N1849);
and AND2 (N3902, N3877, N2901);
buf BUF1 (N3903, N3895);
xor XOR2 (N3904, N3903, N2724);
and AND3 (N3905, N3894, N127, N127);
buf BUF1 (N3906, N3893);
buf BUF1 (N3907, N3901);
nor NOR3 (N3908, N3892, N2207, N1263);
xor XOR2 (N3909, N3897, N3096);
and AND3 (N3910, N3880, N1779, N2421);
nand NAND2 (N3911, N3907, N3798);
or OR2 (N3912, N3905, N3494);
buf BUF1 (N3913, N3902);
and AND2 (N3914, N3906, N3506);
and AND2 (N3915, N3910, N366);
and AND3 (N3916, N3898, N2829, N2768);
xor XOR2 (N3917, N3904, N112);
nand NAND2 (N3918, N3909, N2053);
not NOT1 (N3919, N3908);
or OR3 (N3920, N3887, N200, N2511);
and AND3 (N3921, N3912, N2983, N2314);
not NOT1 (N3922, N3911);
buf BUF1 (N3923, N3913);
nand NAND2 (N3924, N3918, N1941);
not NOT1 (N3925, N3919);
nor NOR4 (N3926, N3923, N3063, N1160, N2499);
nor NOR4 (N3927, N3914, N2053, N1196, N2573);
xor XOR2 (N3928, N3926, N3194);
not NOT1 (N3929, N3917);
xor XOR2 (N3930, N3929, N1599);
or OR2 (N3931, N3928, N2032);
not NOT1 (N3932, N3915);
xor XOR2 (N3933, N3930, N3257);
and AND3 (N3934, N3924, N1908, N3503);
nor NOR2 (N3935, N3931, N1690);
xor XOR2 (N3936, N3933, N3183);
nand NAND2 (N3937, N3932, N3804);
not NOT1 (N3938, N3937);
nand NAND2 (N3939, N3936, N1251);
xor XOR2 (N3940, N3934, N3004);
or OR2 (N3941, N3935, N1547);
buf BUF1 (N3942, N3921);
not NOT1 (N3943, N3938);
xor XOR2 (N3944, N3916, N2547);
and AND2 (N3945, N3943, N704);
nand NAND2 (N3946, N3940, N887);
xor XOR2 (N3947, N3939, N2092);
nand NAND3 (N3948, N3925, N3894, N681);
buf BUF1 (N3949, N3922);
buf BUF1 (N3950, N3942);
buf BUF1 (N3951, N3947);
xor XOR2 (N3952, N3949, N1589);
buf BUF1 (N3953, N3952);
xor XOR2 (N3954, N3944, N394);
or OR2 (N3955, N3927, N2503);
nor NOR3 (N3956, N3948, N2340, N2229);
xor XOR2 (N3957, N3956, N3629);
not NOT1 (N3958, N3953);
or OR2 (N3959, N3950, N2707);
nand NAND4 (N3960, N3945, N2741, N1318, N3225);
or OR3 (N3961, N3960, N312, N3625);
nand NAND4 (N3962, N3954, N1265, N3935, N840);
nand NAND4 (N3963, N3962, N1403, N1657, N1401);
xor XOR2 (N3964, N3951, N1170);
nor NOR2 (N3965, N3955, N667);
and AND4 (N3966, N3957, N1584, N806, N2319);
or OR4 (N3967, N3965, N3324, N1091, N1913);
or OR3 (N3968, N3964, N1361, N55);
xor XOR2 (N3969, N3920, N2866);
nand NAND4 (N3970, N3963, N920, N3359, N2023);
or OR3 (N3971, N3961, N3712, N1883);
xor XOR2 (N3972, N3967, N2729);
nand NAND2 (N3973, N3946, N2325);
nor NOR4 (N3974, N3973, N1177, N1768, N105);
xor XOR2 (N3975, N3969, N3546);
or OR3 (N3976, N3941, N375, N346);
or OR2 (N3977, N3959, N949);
buf BUF1 (N3978, N3958);
or OR2 (N3979, N3971, N3117);
and AND3 (N3980, N3979, N1142, N2156);
nand NAND3 (N3981, N3974, N1361, N3163);
or OR3 (N3982, N3966, N3152, N3424);
buf BUF1 (N3983, N3975);
and AND2 (N3984, N3981, N3285);
buf BUF1 (N3985, N3980);
nand NAND4 (N3986, N3970, N3904, N3697, N1748);
nand NAND2 (N3987, N3985, N3053);
nor NOR3 (N3988, N3983, N1060, N2297);
not NOT1 (N3989, N3968);
nor NOR4 (N3990, N3987, N490, N3722, N3835);
and AND2 (N3991, N3972, N1490);
or OR4 (N3992, N3986, N878, N488, N1047);
buf BUF1 (N3993, N3977);
or OR4 (N3994, N3990, N492, N1285, N94);
or OR3 (N3995, N3982, N2417, N3370);
nand NAND3 (N3996, N3992, N3050, N3919);
not NOT1 (N3997, N3978);
not NOT1 (N3998, N3995);
nor NOR4 (N3999, N3997, N3565, N1606, N2097);
buf BUF1 (N4000, N3991);
or OR2 (N4001, N3996, N3695);
xor XOR2 (N4002, N3993, N877);
nor NOR2 (N4003, N3989, N2871);
not NOT1 (N4004, N4000);
and AND2 (N4005, N4003, N2162);
xor XOR2 (N4006, N3999, N3500);
not NOT1 (N4007, N4006);
buf BUF1 (N4008, N3984);
xor XOR2 (N4009, N4004, N3235);
buf BUF1 (N4010, N3976);
xor XOR2 (N4011, N4001, N2964);
nand NAND2 (N4012, N4010, N1753);
xor XOR2 (N4013, N4008, N1331);
nor NOR2 (N4014, N4005, N1819);
not NOT1 (N4015, N3994);
xor XOR2 (N4016, N4011, N3620);
nor NOR4 (N4017, N3988, N2643, N3385, N1530);
nor NOR4 (N4018, N4012, N737, N585, N504);
xor XOR2 (N4019, N4015, N3307);
buf BUF1 (N4020, N4009);
nand NAND4 (N4021, N4020, N1681, N338, N1712);
nand NAND4 (N4022, N4019, N3406, N2385, N293);
or OR2 (N4023, N4002, N3156);
endmodule