// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17;

output N4008,N4016,N4014,N4012,N4013,N4005,N3989,N3991,N4007,N4017;

buf BUF1 (N18, N2);
not NOT1 (N19, N12);
nor NOR4 (N20, N10, N7, N8, N6);
not NOT1 (N21, N4);
not NOT1 (N22, N10);
nand NAND2 (N23, N22, N21);
nand NAND2 (N24, N23, N23);
or OR2 (N25, N13, N17);
buf BUF1 (N26, N23);
not NOT1 (N27, N18);
not NOT1 (N28, N23);
or OR4 (N29, N14, N11, N1, N18);
buf BUF1 (N30, N28);
xor XOR2 (N31, N26, N8);
nand NAND2 (N32, N30, N31);
and AND2 (N33, N21, N29);
not NOT1 (N34, N18);
nand NAND3 (N35, N10, N8, N22);
buf BUF1 (N36, N18);
not NOT1 (N37, N36);
buf BUF1 (N38, N35);
or OR4 (N39, N34, N11, N20, N32);
xor XOR2 (N40, N31, N3);
and AND2 (N41, N21, N5);
buf BUF1 (N42, N37);
xor XOR2 (N43, N19, N13);
buf BUF1 (N44, N40);
or OR4 (N45, N38, N6, N6, N12);
not NOT1 (N46, N24);
nand NAND3 (N47, N33, N12, N45);
xor XOR2 (N48, N9, N38);
not NOT1 (N49, N42);
or OR3 (N50, N49, N11, N35);
not NOT1 (N51, N25);
or OR4 (N52, N51, N5, N8, N51);
xor XOR2 (N53, N44, N29);
nor NOR4 (N54, N43, N28, N39, N40);
xor XOR2 (N55, N35, N19);
buf BUF1 (N56, N52);
or OR3 (N57, N53, N5, N31);
nor NOR3 (N58, N48, N31, N5);
or OR2 (N59, N56, N5);
and AND3 (N60, N47, N11, N39);
xor XOR2 (N61, N55, N12);
not NOT1 (N62, N41);
not NOT1 (N63, N57);
nand NAND3 (N64, N27, N3, N19);
nor NOR2 (N65, N61, N60);
or OR3 (N66, N17, N22, N20);
not NOT1 (N67, N62);
xor XOR2 (N68, N63, N50);
nand NAND4 (N69, N14, N42, N26, N25);
buf BUF1 (N70, N65);
xor XOR2 (N71, N70, N19);
not NOT1 (N72, N58);
nor NOR4 (N73, N46, N36, N47, N1);
or OR3 (N74, N69, N58, N73);
buf BUF1 (N75, N70);
not NOT1 (N76, N64);
nand NAND4 (N77, N71, N50, N17, N38);
buf BUF1 (N78, N66);
nand NAND4 (N79, N74, N33, N11, N36);
or OR2 (N80, N78, N58);
nand NAND3 (N81, N80, N18, N18);
nand NAND3 (N82, N75, N2, N22);
nand NAND2 (N83, N79, N11);
nor NOR4 (N84, N81, N71, N58, N40);
nand NAND4 (N85, N82, N41, N8, N46);
nor NOR4 (N86, N76, N31, N79, N82);
buf BUF1 (N87, N77);
nand NAND2 (N88, N59, N47);
or OR3 (N89, N68, N65, N88);
nand NAND4 (N90, N75, N62, N81, N44);
not NOT1 (N91, N87);
and AND3 (N92, N67, N78, N49);
nor NOR3 (N93, N83, N84, N47);
not NOT1 (N94, N57);
nor NOR4 (N95, N85, N12, N52, N58);
not NOT1 (N96, N93);
and AND3 (N97, N86, N42, N91);
and AND3 (N98, N28, N55, N64);
not NOT1 (N99, N90);
buf BUF1 (N100, N89);
nand NAND4 (N101, N92, N32, N24, N77);
nor NOR2 (N102, N97, N40);
nand NAND3 (N103, N96, N22, N39);
not NOT1 (N104, N102);
nand NAND3 (N105, N103, N55, N12);
not NOT1 (N106, N99);
buf BUF1 (N107, N104);
xor XOR2 (N108, N106, N14);
xor XOR2 (N109, N107, N53);
nor NOR4 (N110, N101, N100, N49, N109);
nand NAND4 (N111, N26, N52, N38, N29);
not NOT1 (N112, N8);
not NOT1 (N113, N94);
nand NAND2 (N114, N110, N81);
buf BUF1 (N115, N54);
nor NOR3 (N116, N113, N1, N50);
or OR4 (N117, N116, N72, N75, N20);
xor XOR2 (N118, N56, N86);
not NOT1 (N119, N117);
or OR4 (N120, N114, N8, N54, N84);
or OR4 (N121, N112, N116, N81, N39);
and AND2 (N122, N119, N94);
not NOT1 (N123, N95);
or OR2 (N124, N108, N6);
nand NAND2 (N125, N122, N16);
buf BUF1 (N126, N118);
and AND4 (N127, N124, N19, N24, N58);
or OR2 (N128, N121, N107);
or OR4 (N129, N126, N95, N3, N3);
buf BUF1 (N130, N115);
buf BUF1 (N131, N111);
and AND4 (N132, N130, N23, N96, N7);
buf BUF1 (N133, N131);
xor XOR2 (N134, N127, N67);
nor NOR3 (N135, N98, N33, N103);
or OR4 (N136, N125, N74, N99, N78);
buf BUF1 (N137, N123);
not NOT1 (N138, N133);
buf BUF1 (N139, N129);
buf BUF1 (N140, N135);
buf BUF1 (N141, N140);
nor NOR3 (N142, N136, N6, N33);
or OR4 (N143, N120, N6, N34, N121);
xor XOR2 (N144, N128, N112);
and AND3 (N145, N143, N135, N112);
buf BUF1 (N146, N137);
xor XOR2 (N147, N142, N109);
xor XOR2 (N148, N145, N34);
not NOT1 (N149, N139);
nand NAND3 (N150, N147, N146, N69);
nand NAND2 (N151, N98, N6);
nor NOR2 (N152, N132, N49);
buf BUF1 (N153, N138);
nand NAND2 (N154, N151, N110);
buf BUF1 (N155, N141);
buf BUF1 (N156, N148);
nand NAND4 (N157, N149, N116, N32, N71);
not NOT1 (N158, N157);
xor XOR2 (N159, N156, N158);
nand NAND4 (N160, N96, N4, N118, N128);
not NOT1 (N161, N150);
nor NOR2 (N162, N105, N148);
nor NOR4 (N163, N154, N83, N10, N144);
or OR2 (N164, N8, N107);
or OR3 (N165, N164, N21, N73);
nand NAND2 (N166, N163, N29);
or OR3 (N167, N162, N140, N100);
nand NAND4 (N168, N166, N21, N15, N150);
xor XOR2 (N169, N168, N67);
nor NOR2 (N170, N153, N64);
not NOT1 (N171, N152);
xor XOR2 (N172, N134, N25);
nand NAND4 (N173, N172, N129, N155, N96);
and AND2 (N174, N54, N146);
not NOT1 (N175, N170);
and AND4 (N176, N159, N30, N99, N85);
xor XOR2 (N177, N167, N60);
not NOT1 (N178, N173);
or OR4 (N179, N178, N165, N146, N62);
nand NAND3 (N180, N55, N135, N26);
nor NOR2 (N181, N177, N120);
and AND3 (N182, N160, N50, N4);
nand NAND4 (N183, N161, N101, N148, N163);
not NOT1 (N184, N181);
buf BUF1 (N185, N184);
nand NAND4 (N186, N183, N127, N147, N153);
nor NOR2 (N187, N185, N162);
nor NOR3 (N188, N180, N133, N1);
or OR2 (N189, N182, N36);
or OR2 (N190, N187, N141);
not NOT1 (N191, N176);
not NOT1 (N192, N186);
nor NOR3 (N193, N190, N56, N147);
not NOT1 (N194, N192);
buf BUF1 (N195, N171);
and AND2 (N196, N191, N15);
not NOT1 (N197, N194);
buf BUF1 (N198, N179);
not NOT1 (N199, N193);
not NOT1 (N200, N189);
nor NOR2 (N201, N175, N54);
nor NOR2 (N202, N174, N172);
buf BUF1 (N203, N202);
and AND4 (N204, N188, N125, N171, N144);
nor NOR4 (N205, N196, N63, N48, N111);
not NOT1 (N206, N200);
and AND3 (N207, N197, N25, N56);
buf BUF1 (N208, N169);
not NOT1 (N209, N208);
nor NOR2 (N210, N207, N152);
nand NAND2 (N211, N209, N61);
buf BUF1 (N212, N211);
xor XOR2 (N213, N198, N176);
buf BUF1 (N214, N206);
or OR2 (N215, N195, N70);
nand NAND4 (N216, N213, N102, N196, N68);
and AND2 (N217, N212, N112);
nand NAND2 (N218, N216, N35);
and AND4 (N219, N218, N52, N54, N14);
xor XOR2 (N220, N203, N130);
not NOT1 (N221, N199);
buf BUF1 (N222, N214);
and AND3 (N223, N215, N174, N1);
buf BUF1 (N224, N210);
not NOT1 (N225, N224);
nand NAND2 (N226, N222, N207);
or OR2 (N227, N223, N223);
buf BUF1 (N228, N204);
nand NAND4 (N229, N226, N126, N186, N165);
nor NOR3 (N230, N228, N150, N215);
or OR3 (N231, N205, N126, N79);
buf BUF1 (N232, N227);
not NOT1 (N233, N225);
xor XOR2 (N234, N229, N198);
nor NOR2 (N235, N201, N144);
or OR3 (N236, N234, N1, N230);
and AND4 (N237, N146, N234, N192, N54);
or OR3 (N238, N219, N231, N184);
or OR4 (N239, N185, N4, N70, N41);
not NOT1 (N240, N232);
xor XOR2 (N241, N237, N151);
buf BUF1 (N242, N233);
xor XOR2 (N243, N242, N43);
and AND2 (N244, N241, N199);
buf BUF1 (N245, N243);
not NOT1 (N246, N240);
or OR2 (N247, N246, N160);
and AND4 (N248, N220, N64, N85, N134);
nand NAND4 (N249, N217, N190, N126, N35);
and AND4 (N250, N248, N226, N222, N137);
buf BUF1 (N251, N235);
and AND2 (N252, N239, N197);
nand NAND2 (N253, N249, N77);
buf BUF1 (N254, N236);
or OR4 (N255, N221, N76, N10, N64);
or OR3 (N256, N247, N238, N232);
and AND3 (N257, N211, N202, N58);
nor NOR3 (N258, N250, N189, N21);
or OR3 (N259, N254, N96, N50);
and AND3 (N260, N252, N233, N177);
not NOT1 (N261, N245);
nand NAND4 (N262, N260, N39, N44, N232);
buf BUF1 (N263, N251);
not NOT1 (N264, N259);
nand NAND2 (N265, N262, N156);
and AND2 (N266, N244, N74);
nand NAND4 (N267, N263, N125, N226, N176);
or OR3 (N268, N264, N81, N182);
not NOT1 (N269, N266);
not NOT1 (N270, N257);
nand NAND3 (N271, N268, N107, N58);
or OR3 (N272, N261, N56, N85);
nand NAND2 (N273, N255, N189);
nand NAND2 (N274, N273, N169);
not NOT1 (N275, N267);
and AND4 (N276, N274, N88, N75, N259);
nand NAND3 (N277, N253, N155, N166);
xor XOR2 (N278, N256, N72);
or OR4 (N279, N277, N208, N102, N163);
and AND4 (N280, N258, N112, N15, N67);
or OR3 (N281, N272, N263, N33);
nand NAND3 (N282, N276, N251, N90);
nand NAND3 (N283, N269, N97, N116);
nor NOR3 (N284, N271, N196, N63);
buf BUF1 (N285, N270);
not NOT1 (N286, N280);
or OR2 (N287, N279, N114);
nor NOR4 (N288, N287, N181, N42, N65);
xor XOR2 (N289, N275, N284);
not NOT1 (N290, N87);
nor NOR3 (N291, N288, N35, N152);
nand NAND4 (N292, N283, N177, N166, N160);
not NOT1 (N293, N278);
or OR4 (N294, N286, N102, N161, N118);
nand NAND3 (N295, N265, N154, N17);
not NOT1 (N296, N282);
not NOT1 (N297, N281);
nand NAND4 (N298, N290, N80, N73, N71);
not NOT1 (N299, N294);
xor XOR2 (N300, N293, N261);
nand NAND2 (N301, N292, N141);
xor XOR2 (N302, N291, N214);
nor NOR3 (N303, N300, N223, N89);
xor XOR2 (N304, N297, N163);
not NOT1 (N305, N295);
or OR2 (N306, N298, N203);
nand NAND3 (N307, N302, N150, N20);
nor NOR4 (N308, N285, N259, N60, N119);
nand NAND4 (N309, N301, N222, N23, N23);
not NOT1 (N310, N303);
buf BUF1 (N311, N310);
not NOT1 (N312, N311);
xor XOR2 (N313, N296, N123);
or OR3 (N314, N299, N120, N75);
and AND4 (N315, N312, N165, N35, N40);
nor NOR4 (N316, N306, N239, N12, N258);
xor XOR2 (N317, N316, N47);
nand NAND3 (N318, N289, N248, N114);
and AND3 (N319, N304, N316, N89);
nand NAND3 (N320, N315, N108, N250);
not NOT1 (N321, N305);
or OR3 (N322, N314, N134, N41);
nand NAND3 (N323, N322, N186, N117);
nand NAND2 (N324, N323, N26);
not NOT1 (N325, N309);
xor XOR2 (N326, N318, N158);
xor XOR2 (N327, N324, N247);
buf BUF1 (N328, N308);
not NOT1 (N329, N321);
or OR2 (N330, N329, N276);
and AND4 (N331, N307, N52, N85, N264);
xor XOR2 (N332, N313, N55);
or OR4 (N333, N331, N72, N65, N267);
and AND2 (N334, N328, N309);
and AND3 (N335, N317, N199, N285);
xor XOR2 (N336, N319, N306);
nand NAND2 (N337, N335, N333);
nand NAND3 (N338, N170, N19, N213);
nand NAND3 (N339, N332, N116, N198);
buf BUF1 (N340, N338);
nand NAND2 (N341, N326, N35);
not NOT1 (N342, N341);
buf BUF1 (N343, N320);
not NOT1 (N344, N330);
or OR3 (N345, N343, N273, N246);
buf BUF1 (N346, N342);
buf BUF1 (N347, N325);
or OR2 (N348, N347, N17);
or OR4 (N349, N336, N221, N314, N316);
xor XOR2 (N350, N340, N145);
xor XOR2 (N351, N346, N280);
buf BUF1 (N352, N327);
or OR2 (N353, N348, N203);
nor NOR4 (N354, N339, N332, N148, N173);
not NOT1 (N355, N334);
nand NAND3 (N356, N350, N77, N124);
and AND4 (N357, N355, N229, N285, N30);
nor NOR3 (N358, N354, N244, N247);
or OR4 (N359, N357, N87, N10, N87);
and AND4 (N360, N337, N324, N261, N106);
nand NAND4 (N361, N351, N7, N144, N68);
buf BUF1 (N362, N345);
nand NAND3 (N363, N344, N269, N254);
nor NOR4 (N364, N352, N109, N51, N24);
and AND3 (N365, N359, N61, N268);
xor XOR2 (N366, N358, N86);
or OR2 (N367, N364, N16);
or OR2 (N368, N362, N267);
nand NAND3 (N369, N360, N239, N332);
nor NOR4 (N370, N369, N177, N266, N32);
xor XOR2 (N371, N365, N45);
nor NOR3 (N372, N371, N11, N50);
xor XOR2 (N373, N366, N67);
nor NOR4 (N374, N373, N12, N208, N171);
xor XOR2 (N375, N368, N205);
buf BUF1 (N376, N370);
or OR2 (N377, N363, N24);
nand NAND2 (N378, N356, N251);
buf BUF1 (N379, N377);
buf BUF1 (N380, N372);
nor NOR2 (N381, N376, N180);
and AND4 (N382, N367, N155, N159, N292);
nand NAND4 (N383, N349, N50, N19, N237);
or OR2 (N384, N381, N25);
or OR2 (N385, N374, N226);
and AND2 (N386, N380, N236);
buf BUF1 (N387, N378);
buf BUF1 (N388, N361);
or OR4 (N389, N379, N285, N336, N3);
or OR2 (N390, N375, N344);
nor NOR4 (N391, N382, N167, N325, N289);
not NOT1 (N392, N390);
nor NOR2 (N393, N385, N16);
nor NOR3 (N394, N388, N357, N49);
or OR4 (N395, N387, N217, N76, N320);
nand NAND3 (N396, N384, N390, N109);
not NOT1 (N397, N394);
xor XOR2 (N398, N395, N167);
or OR2 (N399, N397, N358);
xor XOR2 (N400, N396, N161);
and AND4 (N401, N389, N6, N17, N21);
nand NAND4 (N402, N401, N393, N71, N80);
not NOT1 (N403, N392);
buf BUF1 (N404, N391);
nand NAND2 (N405, N3, N315);
not NOT1 (N406, N402);
nand NAND2 (N407, N383, N324);
buf BUF1 (N408, N403);
and AND4 (N409, N404, N294, N41, N164);
xor XOR2 (N410, N409, N231);
nand NAND4 (N411, N353, N244, N209, N234);
buf BUF1 (N412, N405);
or OR3 (N413, N399, N167, N160);
buf BUF1 (N414, N410);
and AND2 (N415, N413, N366);
nor NOR2 (N416, N407, N208);
xor XOR2 (N417, N412, N288);
xor XOR2 (N418, N414, N411);
xor XOR2 (N419, N220, N124);
buf BUF1 (N420, N415);
and AND2 (N421, N419, N54);
nand NAND2 (N422, N417, N35);
buf BUF1 (N423, N418);
buf BUF1 (N424, N400);
xor XOR2 (N425, N406, N394);
xor XOR2 (N426, N420, N251);
nor NOR4 (N427, N425, N161, N344, N148);
and AND2 (N428, N422, N317);
buf BUF1 (N429, N426);
or OR2 (N430, N429, N47);
xor XOR2 (N431, N408, N261);
nand NAND4 (N432, N421, N420, N171, N317);
nand NAND2 (N433, N427, N193);
nand NAND4 (N434, N423, N49, N94, N298);
and AND3 (N435, N424, N316, N274);
buf BUF1 (N436, N434);
buf BUF1 (N437, N398);
not NOT1 (N438, N416);
xor XOR2 (N439, N430, N153);
nor NOR3 (N440, N431, N137, N397);
or OR4 (N441, N433, N182, N384, N260);
buf BUF1 (N442, N439);
and AND4 (N443, N441, N180, N372, N206);
nand NAND2 (N444, N435, N137);
buf BUF1 (N445, N437);
or OR4 (N446, N443, N13, N426, N290);
buf BUF1 (N447, N445);
nor NOR3 (N448, N386, N44, N447);
not NOT1 (N449, N396);
nand NAND2 (N450, N428, N148);
xor XOR2 (N451, N450, N139);
nand NAND4 (N452, N446, N207, N441, N302);
buf BUF1 (N453, N442);
or OR4 (N454, N436, N318, N202, N131);
not NOT1 (N455, N432);
nor NOR2 (N456, N440, N118);
buf BUF1 (N457, N449);
xor XOR2 (N458, N456, N251);
nand NAND2 (N459, N455, N259);
xor XOR2 (N460, N451, N266);
nand NAND3 (N461, N454, N392, N401);
xor XOR2 (N462, N459, N244);
not NOT1 (N463, N457);
not NOT1 (N464, N460);
xor XOR2 (N465, N463, N386);
buf BUF1 (N466, N464);
nor NOR3 (N467, N466, N406, N326);
buf BUF1 (N468, N444);
or OR2 (N469, N438, N284);
xor XOR2 (N470, N462, N442);
xor XOR2 (N471, N448, N93);
not NOT1 (N472, N469);
nor NOR4 (N473, N461, N57, N259, N468);
and AND4 (N474, N170, N192, N388, N366);
nor NOR4 (N475, N465, N197, N155, N66);
nor NOR3 (N476, N470, N98, N144);
buf BUF1 (N477, N452);
nand NAND3 (N478, N474, N304, N298);
and AND2 (N479, N477, N73);
nand NAND4 (N480, N475, N473, N252, N281);
xor XOR2 (N481, N19, N480);
nand NAND2 (N482, N82, N125);
buf BUF1 (N483, N479);
xor XOR2 (N484, N453, N187);
not NOT1 (N485, N476);
nand NAND3 (N486, N458, N143, N446);
and AND4 (N487, N486, N360, N111, N271);
buf BUF1 (N488, N467);
or OR2 (N489, N485, N152);
not NOT1 (N490, N489);
or OR3 (N491, N490, N11, N120);
not NOT1 (N492, N491);
or OR2 (N493, N487, N127);
or OR2 (N494, N493, N458);
buf BUF1 (N495, N482);
nor NOR4 (N496, N471, N413, N24, N52);
not NOT1 (N497, N496);
not NOT1 (N498, N472);
buf BUF1 (N499, N478);
and AND4 (N500, N499, N40, N6, N489);
and AND4 (N501, N497, N379, N428, N425);
not NOT1 (N502, N500);
buf BUF1 (N503, N501);
nand NAND2 (N504, N481, N483);
nor NOR4 (N505, N77, N58, N390, N488);
not NOT1 (N506, N224);
or OR2 (N507, N494, N489);
not NOT1 (N508, N495);
not NOT1 (N509, N505);
nand NAND3 (N510, N503, N136, N320);
nor NOR4 (N511, N502, N467, N414, N134);
and AND2 (N512, N484, N503);
xor XOR2 (N513, N510, N464);
not NOT1 (N514, N509);
or OR4 (N515, N492, N277, N510, N243);
buf BUF1 (N516, N512);
and AND3 (N517, N498, N245, N228);
buf BUF1 (N518, N513);
not NOT1 (N519, N515);
nor NOR4 (N520, N511, N473, N23, N266);
or OR2 (N521, N517, N141);
nand NAND4 (N522, N504, N507, N295, N409);
or OR4 (N523, N175, N1, N179, N88);
nor NOR2 (N524, N518, N179);
not NOT1 (N525, N523);
or OR4 (N526, N514, N182, N506, N5);
nor NOR4 (N527, N331, N290, N268, N87);
and AND2 (N528, N516, N343);
or OR3 (N529, N520, N60, N319);
or OR3 (N530, N528, N107, N118);
or OR2 (N531, N508, N393);
buf BUF1 (N532, N526);
xor XOR2 (N533, N532, N347);
or OR3 (N534, N527, N371, N246);
or OR2 (N535, N529, N350);
or OR2 (N536, N535, N314);
or OR4 (N537, N534, N372, N334, N261);
xor XOR2 (N538, N521, N223);
xor XOR2 (N539, N531, N410);
not NOT1 (N540, N522);
xor XOR2 (N541, N536, N47);
or OR4 (N542, N519, N10, N210, N397);
nand NAND4 (N543, N540, N10, N68, N25);
not NOT1 (N544, N524);
not NOT1 (N545, N538);
xor XOR2 (N546, N525, N192);
buf BUF1 (N547, N541);
nand NAND4 (N548, N543, N262, N153, N416);
nand NAND4 (N549, N546, N439, N89, N396);
xor XOR2 (N550, N533, N540);
not NOT1 (N551, N545);
or OR3 (N552, N537, N230, N224);
nand NAND3 (N553, N539, N309, N288);
or OR2 (N554, N544, N242);
or OR4 (N555, N550, N37, N441, N343);
or OR4 (N556, N547, N400, N136, N1);
not NOT1 (N557, N548);
or OR3 (N558, N554, N28, N461);
nand NAND2 (N559, N552, N264);
and AND4 (N560, N542, N174, N71, N195);
xor XOR2 (N561, N558, N187);
or OR3 (N562, N557, N257, N163);
nand NAND4 (N563, N560, N178, N251, N304);
xor XOR2 (N564, N563, N258);
or OR2 (N565, N549, N2);
and AND4 (N566, N553, N526, N180, N25);
nand NAND3 (N567, N564, N122, N327);
and AND2 (N568, N561, N232);
or OR4 (N569, N555, N53, N222, N515);
and AND2 (N570, N551, N245);
or OR3 (N571, N567, N373, N463);
not NOT1 (N572, N571);
and AND3 (N573, N562, N234, N119);
nand NAND4 (N574, N566, N220, N409, N329);
not NOT1 (N575, N570);
or OR3 (N576, N530, N424, N25);
xor XOR2 (N577, N575, N77);
buf BUF1 (N578, N574);
buf BUF1 (N579, N576);
xor XOR2 (N580, N572, N477);
and AND4 (N581, N559, N485, N305, N65);
or OR4 (N582, N577, N105, N98, N33);
buf BUF1 (N583, N582);
or OR3 (N584, N579, N261, N281);
xor XOR2 (N585, N573, N44);
or OR3 (N586, N585, N488, N27);
nor NOR3 (N587, N565, N451, N195);
or OR4 (N588, N556, N146, N380, N273);
nand NAND4 (N589, N583, N217, N366, N158);
nor NOR2 (N590, N588, N503);
not NOT1 (N591, N581);
or OR2 (N592, N578, N400);
buf BUF1 (N593, N592);
not NOT1 (N594, N587);
nand NAND4 (N595, N591, N382, N137, N251);
or OR2 (N596, N595, N378);
or OR2 (N597, N596, N355);
and AND2 (N598, N580, N284);
not NOT1 (N599, N594);
nand NAND2 (N600, N589, N500);
buf BUF1 (N601, N584);
and AND2 (N602, N601, N207);
buf BUF1 (N603, N590);
and AND3 (N604, N568, N591, N12);
xor XOR2 (N605, N569, N284);
nor NOR2 (N606, N604, N76);
xor XOR2 (N607, N586, N344);
nor NOR4 (N608, N606, N588, N517, N423);
nand NAND2 (N609, N602, N493);
not NOT1 (N610, N593);
buf BUF1 (N611, N599);
buf BUF1 (N612, N611);
not NOT1 (N613, N603);
xor XOR2 (N614, N612, N230);
buf BUF1 (N615, N600);
and AND2 (N616, N597, N443);
and AND4 (N617, N608, N65, N495, N462);
xor XOR2 (N618, N613, N278);
nand NAND4 (N619, N607, N519, N421, N482);
nor NOR2 (N620, N614, N302);
nand NAND2 (N621, N609, N526);
nor NOR4 (N622, N618, N471, N297, N128);
xor XOR2 (N623, N605, N601);
not NOT1 (N624, N616);
or OR2 (N625, N615, N311);
or OR2 (N626, N620, N163);
nor NOR3 (N627, N626, N133, N520);
nand NAND3 (N628, N622, N391, N270);
buf BUF1 (N629, N621);
not NOT1 (N630, N628);
or OR2 (N631, N598, N288);
buf BUF1 (N632, N610);
buf BUF1 (N633, N623);
nor NOR3 (N634, N627, N55, N447);
buf BUF1 (N635, N634);
nand NAND4 (N636, N617, N541, N517, N315);
nand NAND4 (N637, N629, N160, N431, N206);
nor NOR4 (N638, N624, N165, N333, N11);
and AND4 (N639, N635, N478, N377, N280);
buf BUF1 (N640, N637);
nand NAND3 (N641, N639, N421, N8);
nor NOR4 (N642, N638, N22, N149, N188);
buf BUF1 (N643, N636);
and AND4 (N644, N632, N373, N139, N599);
or OR3 (N645, N631, N378, N585);
and AND4 (N646, N645, N271, N554, N123);
nor NOR2 (N647, N642, N160);
buf BUF1 (N648, N647);
buf BUF1 (N649, N641);
nand NAND4 (N650, N640, N263, N570, N308);
xor XOR2 (N651, N648, N548);
or OR4 (N652, N651, N339, N457, N481);
xor XOR2 (N653, N650, N620);
or OR4 (N654, N643, N519, N130, N184);
or OR4 (N655, N654, N497, N624, N463);
nor NOR4 (N656, N630, N318, N321, N480);
xor XOR2 (N657, N656, N511);
not NOT1 (N658, N633);
nand NAND2 (N659, N619, N103);
not NOT1 (N660, N652);
or OR2 (N661, N658, N161);
buf BUF1 (N662, N649);
nand NAND3 (N663, N653, N498, N358);
not NOT1 (N664, N663);
and AND3 (N665, N625, N145, N663);
not NOT1 (N666, N657);
buf BUF1 (N667, N665);
nor NOR4 (N668, N644, N435, N455, N619);
nand NAND4 (N669, N661, N278, N51, N324);
and AND3 (N670, N655, N441, N606);
buf BUF1 (N671, N668);
not NOT1 (N672, N667);
nand NAND2 (N673, N659, N55);
not NOT1 (N674, N646);
and AND3 (N675, N662, N236, N557);
buf BUF1 (N676, N664);
nor NOR2 (N677, N670, N162);
nand NAND2 (N678, N672, N462);
or OR3 (N679, N674, N330, N324);
nand NAND2 (N680, N671, N634);
xor XOR2 (N681, N680, N363);
and AND2 (N682, N681, N201);
or OR3 (N683, N669, N540, N479);
xor XOR2 (N684, N673, N255);
or OR3 (N685, N684, N585, N32);
xor XOR2 (N686, N666, N526);
nor NOR3 (N687, N678, N351, N50);
buf BUF1 (N688, N675);
or OR2 (N689, N688, N453);
nand NAND3 (N690, N689, N477, N132);
and AND3 (N691, N686, N280, N620);
nand NAND3 (N692, N660, N427, N68);
nand NAND2 (N693, N691, N489);
nand NAND4 (N694, N677, N77, N52, N582);
not NOT1 (N695, N682);
or OR4 (N696, N693, N314, N622, N567);
nand NAND4 (N697, N676, N516, N577, N572);
buf BUF1 (N698, N696);
nor NOR3 (N699, N679, N522, N674);
and AND2 (N700, N695, N143);
xor XOR2 (N701, N694, N59);
buf BUF1 (N702, N685);
and AND2 (N703, N690, N496);
and AND2 (N704, N699, N559);
not NOT1 (N705, N701);
not NOT1 (N706, N697);
or OR2 (N707, N706, N544);
or OR4 (N708, N683, N385, N704, N475);
or OR4 (N709, N196, N707, N580, N160);
nand NAND2 (N710, N476, N100);
not NOT1 (N711, N710);
not NOT1 (N712, N698);
not NOT1 (N713, N712);
nor NOR2 (N714, N708, N78);
or OR3 (N715, N687, N314, N376);
and AND4 (N716, N692, N633, N698, N489);
nor NOR4 (N717, N713, N261, N415, N79);
not NOT1 (N718, N715);
buf BUF1 (N719, N703);
nand NAND4 (N720, N700, N679, N484, N399);
not NOT1 (N721, N702);
nand NAND2 (N722, N711, N600);
buf BUF1 (N723, N721);
and AND4 (N724, N719, N365, N652, N177);
buf BUF1 (N725, N724);
nor NOR3 (N726, N716, N511, N533);
buf BUF1 (N727, N705);
nor NOR2 (N728, N714, N251);
or OR4 (N729, N718, N633, N591, N318);
or OR3 (N730, N728, N498, N207);
nand NAND3 (N731, N722, N537, N609);
or OR3 (N732, N723, N637, N611);
or OR2 (N733, N727, N295);
buf BUF1 (N734, N726);
buf BUF1 (N735, N730);
not NOT1 (N736, N734);
or OR3 (N737, N735, N261, N521);
or OR3 (N738, N731, N465, N574);
not NOT1 (N739, N732);
xor XOR2 (N740, N737, N577);
buf BUF1 (N741, N733);
buf BUF1 (N742, N741);
nand NAND3 (N743, N717, N706, N197);
buf BUF1 (N744, N739);
buf BUF1 (N745, N738);
buf BUF1 (N746, N740);
or OR4 (N747, N746, N682, N37, N481);
nor NOR3 (N748, N744, N519, N715);
nand NAND3 (N749, N742, N95, N375);
nor NOR4 (N750, N709, N718, N468, N667);
and AND4 (N751, N720, N743, N236, N737);
or OR3 (N752, N371, N620, N299);
nand NAND3 (N753, N747, N305, N603);
and AND3 (N754, N753, N285, N537);
buf BUF1 (N755, N748);
and AND2 (N756, N736, N276);
or OR2 (N757, N745, N614);
buf BUF1 (N758, N725);
nand NAND3 (N759, N729, N129, N757);
not NOT1 (N760, N100);
or OR3 (N761, N752, N520, N202);
xor XOR2 (N762, N749, N67);
nand NAND2 (N763, N756, N320);
nor NOR4 (N764, N760, N431, N473, N116);
nand NAND2 (N765, N763, N367);
or OR2 (N766, N755, N94);
nand NAND3 (N767, N759, N532, N672);
buf BUF1 (N768, N762);
xor XOR2 (N769, N761, N330);
and AND4 (N770, N765, N234, N132, N229);
and AND3 (N771, N750, N374, N686);
or OR2 (N772, N767, N719);
xor XOR2 (N773, N772, N652);
not NOT1 (N774, N758);
and AND3 (N775, N770, N493, N23);
not NOT1 (N776, N751);
xor XOR2 (N777, N766, N15);
xor XOR2 (N778, N773, N5);
and AND2 (N779, N769, N590);
nor NOR4 (N780, N768, N125, N499, N73);
nor NOR3 (N781, N775, N714, N646);
nor NOR2 (N782, N777, N569);
nor NOR2 (N783, N781, N761);
xor XOR2 (N784, N776, N608);
not NOT1 (N785, N771);
xor XOR2 (N786, N778, N39);
buf BUF1 (N787, N783);
xor XOR2 (N788, N774, N445);
buf BUF1 (N789, N782);
and AND4 (N790, N788, N140, N218, N162);
and AND3 (N791, N789, N129, N148);
nor NOR2 (N792, N780, N321);
and AND3 (N793, N786, N90, N553);
nor NOR4 (N794, N785, N24, N654, N370);
xor XOR2 (N795, N793, N221);
or OR3 (N796, N795, N69, N113);
buf BUF1 (N797, N796);
and AND2 (N798, N784, N640);
nand NAND3 (N799, N787, N585, N196);
nand NAND2 (N800, N779, N188);
nand NAND4 (N801, N754, N83, N420, N600);
xor XOR2 (N802, N794, N745);
xor XOR2 (N803, N802, N735);
nand NAND2 (N804, N764, N304);
or OR3 (N805, N800, N524, N142);
nand NAND3 (N806, N804, N342, N794);
and AND3 (N807, N806, N538, N186);
xor XOR2 (N808, N805, N11);
xor XOR2 (N809, N798, N435);
buf BUF1 (N810, N807);
and AND3 (N811, N799, N606, N254);
not NOT1 (N812, N791);
and AND2 (N813, N812, N4);
nand NAND3 (N814, N797, N483, N796);
nor NOR3 (N815, N813, N501, N391);
not NOT1 (N816, N809);
buf BUF1 (N817, N810);
xor XOR2 (N818, N792, N270);
buf BUF1 (N819, N817);
or OR2 (N820, N815, N317);
not NOT1 (N821, N803);
nor NOR3 (N822, N808, N270, N540);
buf BUF1 (N823, N821);
nand NAND2 (N824, N816, N633);
nand NAND3 (N825, N814, N694, N327);
and AND3 (N826, N818, N716, N655);
or OR4 (N827, N801, N545, N29, N397);
not NOT1 (N828, N811);
xor XOR2 (N829, N824, N392);
nor NOR3 (N830, N823, N121, N303);
not NOT1 (N831, N822);
nand NAND4 (N832, N827, N773, N503, N518);
nor NOR2 (N833, N828, N696);
nand NAND4 (N834, N826, N113, N800, N328);
nand NAND3 (N835, N834, N623, N121);
not NOT1 (N836, N832);
and AND2 (N837, N825, N223);
or OR2 (N838, N833, N808);
nand NAND2 (N839, N838, N23);
buf BUF1 (N840, N819);
nand NAND2 (N841, N831, N56);
nor NOR4 (N842, N830, N582, N2, N283);
or OR2 (N843, N820, N183);
and AND3 (N844, N842, N119, N328);
xor XOR2 (N845, N840, N363);
buf BUF1 (N846, N836);
or OR3 (N847, N829, N92, N784);
buf BUF1 (N848, N846);
buf BUF1 (N849, N839);
and AND4 (N850, N845, N522, N313, N496);
nor NOR3 (N851, N790, N612, N550);
buf BUF1 (N852, N844);
nand NAND4 (N853, N843, N486, N144, N52);
nor NOR3 (N854, N849, N781, N12);
buf BUF1 (N855, N847);
nor NOR3 (N856, N848, N611, N551);
or OR2 (N857, N855, N154);
buf BUF1 (N858, N854);
nor NOR3 (N859, N857, N471, N693);
nor NOR3 (N860, N850, N527, N553);
nand NAND3 (N861, N837, N426, N419);
and AND2 (N862, N841, N726);
nand NAND3 (N863, N835, N426, N650);
and AND4 (N864, N853, N10, N334, N334);
not NOT1 (N865, N858);
not NOT1 (N866, N865);
nand NAND3 (N867, N864, N695, N414);
or OR3 (N868, N866, N641, N683);
buf BUF1 (N869, N862);
or OR2 (N870, N859, N834);
xor XOR2 (N871, N868, N113);
nand NAND3 (N872, N856, N502, N854);
not NOT1 (N873, N872);
nand NAND3 (N874, N867, N384, N831);
or OR3 (N875, N860, N525, N71);
xor XOR2 (N876, N874, N37);
or OR2 (N877, N873, N318);
nand NAND4 (N878, N870, N644, N839, N805);
xor XOR2 (N879, N851, N557);
xor XOR2 (N880, N875, N52);
nand NAND2 (N881, N876, N248);
nand NAND3 (N882, N871, N633, N322);
or OR4 (N883, N861, N37, N452, N628);
or OR2 (N884, N852, N11);
buf BUF1 (N885, N880);
nand NAND2 (N886, N884, N507);
nor NOR2 (N887, N878, N617);
buf BUF1 (N888, N887);
or OR2 (N889, N886, N834);
and AND4 (N890, N885, N497, N439, N420);
xor XOR2 (N891, N877, N40);
nor NOR2 (N892, N879, N176);
xor XOR2 (N893, N890, N171);
or OR3 (N894, N869, N751, N497);
not NOT1 (N895, N893);
and AND4 (N896, N895, N863, N166, N807);
not NOT1 (N897, N500);
xor XOR2 (N898, N889, N638);
xor XOR2 (N899, N892, N79);
or OR2 (N900, N891, N38);
nor NOR3 (N901, N899, N268, N568);
nand NAND4 (N902, N881, N744, N884, N1);
and AND2 (N903, N902, N566);
buf BUF1 (N904, N901);
and AND4 (N905, N882, N528, N593, N95);
not NOT1 (N906, N896);
and AND2 (N907, N903, N700);
not NOT1 (N908, N907);
not NOT1 (N909, N898);
nor NOR4 (N910, N888, N724, N475, N164);
or OR2 (N911, N910, N814);
xor XOR2 (N912, N906, N737);
not NOT1 (N913, N897);
xor XOR2 (N914, N883, N594);
nand NAND3 (N915, N909, N480, N285);
buf BUF1 (N916, N900);
not NOT1 (N917, N911);
nand NAND2 (N918, N908, N420);
nand NAND2 (N919, N904, N324);
xor XOR2 (N920, N913, N40);
or OR2 (N921, N915, N678);
not NOT1 (N922, N894);
nor NOR2 (N923, N912, N412);
xor XOR2 (N924, N917, N507);
nor NOR2 (N925, N916, N116);
buf BUF1 (N926, N918);
or OR2 (N927, N914, N491);
and AND2 (N928, N919, N420);
nor NOR4 (N929, N927, N680, N821, N637);
nand NAND4 (N930, N929, N652, N395, N290);
and AND2 (N931, N926, N148);
nor NOR4 (N932, N930, N67, N678, N86);
not NOT1 (N933, N923);
or OR4 (N934, N920, N852, N860, N305);
and AND3 (N935, N922, N22, N426);
nand NAND2 (N936, N921, N863);
buf BUF1 (N937, N905);
not NOT1 (N938, N932);
nor NOR4 (N939, N938, N822, N889, N598);
buf BUF1 (N940, N924);
not NOT1 (N941, N940);
nand NAND3 (N942, N933, N622, N635);
nor NOR4 (N943, N931, N736, N861, N463);
or OR2 (N944, N942, N757);
buf BUF1 (N945, N928);
nor NOR4 (N946, N925, N409, N730, N103);
not NOT1 (N947, N941);
not NOT1 (N948, N947);
xor XOR2 (N949, N936, N594);
not NOT1 (N950, N945);
nor NOR2 (N951, N943, N196);
buf BUF1 (N952, N949);
and AND3 (N953, N950, N284, N784);
not NOT1 (N954, N948);
or OR3 (N955, N944, N626, N32);
buf BUF1 (N956, N934);
not NOT1 (N957, N939);
buf BUF1 (N958, N955);
buf BUF1 (N959, N958);
buf BUF1 (N960, N954);
not NOT1 (N961, N937);
nand NAND4 (N962, N953, N799, N37, N259);
buf BUF1 (N963, N959);
nand NAND3 (N964, N963, N273, N363);
xor XOR2 (N965, N951, N521);
nand NAND2 (N966, N961, N229);
not NOT1 (N967, N946);
buf BUF1 (N968, N956);
buf BUF1 (N969, N964);
nor NOR2 (N970, N952, N196);
or OR2 (N971, N935, N474);
nor NOR2 (N972, N967, N807);
buf BUF1 (N973, N970);
or OR4 (N974, N962, N281, N102, N742);
and AND3 (N975, N957, N726, N514);
or OR2 (N976, N974, N363);
nand NAND3 (N977, N971, N654, N641);
or OR2 (N978, N976, N885);
nor NOR2 (N979, N978, N333);
nor NOR3 (N980, N977, N786, N267);
xor XOR2 (N981, N960, N914);
and AND4 (N982, N968, N864, N301, N932);
and AND4 (N983, N982, N365, N205, N710);
or OR3 (N984, N983, N887, N710);
nor NOR2 (N985, N975, N752);
xor XOR2 (N986, N985, N351);
nand NAND4 (N987, N973, N608, N723, N309);
or OR4 (N988, N979, N9, N278, N841);
and AND4 (N989, N986, N710, N722, N124);
buf BUF1 (N990, N981);
xor XOR2 (N991, N988, N493);
nand NAND4 (N992, N989, N235, N329, N948);
and AND2 (N993, N980, N433);
and AND3 (N994, N992, N114, N143);
not NOT1 (N995, N972);
and AND3 (N996, N991, N485, N948);
not NOT1 (N997, N969);
nor NOR3 (N998, N965, N255, N380);
and AND4 (N999, N987, N504, N822, N277);
and AND4 (N1000, N999, N328, N74, N411);
xor XOR2 (N1001, N966, N842);
nor NOR2 (N1002, N998, N860);
buf BUF1 (N1003, N997);
nor NOR4 (N1004, N1002, N445, N507, N224);
and AND2 (N1005, N996, N886);
nand NAND2 (N1006, N994, N401);
nand NAND4 (N1007, N990, N655, N117, N753);
buf BUF1 (N1008, N1003);
buf BUF1 (N1009, N1000);
nor NOR4 (N1010, N1005, N918, N532, N174);
xor XOR2 (N1011, N1006, N629);
and AND2 (N1012, N995, N834);
and AND3 (N1013, N1004, N537, N897);
and AND4 (N1014, N1013, N191, N305, N59);
and AND3 (N1015, N1009, N930, N41);
and AND2 (N1016, N1008, N919);
buf BUF1 (N1017, N1014);
xor XOR2 (N1018, N1011, N369);
buf BUF1 (N1019, N1017);
xor XOR2 (N1020, N1016, N306);
nand NAND2 (N1021, N1020, N912);
xor XOR2 (N1022, N1021, N692);
buf BUF1 (N1023, N1019);
and AND4 (N1024, N1018, N768, N112, N704);
buf BUF1 (N1025, N1007);
not NOT1 (N1026, N1022);
buf BUF1 (N1027, N993);
not NOT1 (N1028, N1012);
or OR4 (N1029, N1026, N109, N546, N878);
or OR4 (N1030, N1010, N1009, N170, N705);
or OR2 (N1031, N1027, N449);
nor NOR4 (N1032, N1015, N217, N208, N300);
nor NOR2 (N1033, N1025, N442);
nor NOR3 (N1034, N1031, N362, N271);
and AND4 (N1035, N1030, N684, N970, N838);
nor NOR3 (N1036, N984, N820, N736);
nor NOR4 (N1037, N1028, N300, N1024, N812);
and AND2 (N1038, N322, N339);
not NOT1 (N1039, N1023);
nand NAND2 (N1040, N1038, N702);
xor XOR2 (N1041, N1037, N622);
nor NOR3 (N1042, N1032, N637, N386);
or OR4 (N1043, N1036, N717, N876, N484);
nand NAND2 (N1044, N1041, N37);
or OR3 (N1045, N1034, N800, N717);
or OR4 (N1046, N1001, N178, N47, N771);
nor NOR3 (N1047, N1033, N458, N137);
nor NOR4 (N1048, N1042, N675, N351, N379);
buf BUF1 (N1049, N1046);
not NOT1 (N1050, N1043);
not NOT1 (N1051, N1040);
xor XOR2 (N1052, N1051, N797);
nand NAND4 (N1053, N1050, N802, N605, N204);
not NOT1 (N1054, N1053);
or OR3 (N1055, N1029, N468, N724);
or OR4 (N1056, N1045, N322, N869, N860);
nand NAND2 (N1057, N1054, N535);
buf BUF1 (N1058, N1055);
buf BUF1 (N1059, N1035);
xor XOR2 (N1060, N1049, N144);
or OR3 (N1061, N1052, N427, N974);
xor XOR2 (N1062, N1048, N959);
or OR3 (N1063, N1060, N822, N216);
nor NOR4 (N1064, N1044, N1022, N739, N469);
nand NAND2 (N1065, N1047, N531);
buf BUF1 (N1066, N1065);
buf BUF1 (N1067, N1062);
nand NAND4 (N1068, N1039, N598, N926, N662);
buf BUF1 (N1069, N1061);
nor NOR3 (N1070, N1067, N401, N833);
and AND3 (N1071, N1063, N356, N586);
not NOT1 (N1072, N1058);
and AND3 (N1073, N1059, N867, N776);
nor NOR4 (N1074, N1064, N649, N49, N416);
nor NOR3 (N1075, N1056, N820, N225);
or OR3 (N1076, N1071, N238, N436);
not NOT1 (N1077, N1068);
nor NOR4 (N1078, N1069, N372, N919, N924);
or OR3 (N1079, N1077, N11, N725);
or OR4 (N1080, N1076, N475, N49, N150);
not NOT1 (N1081, N1074);
xor XOR2 (N1082, N1066, N428);
and AND4 (N1083, N1079, N370, N227, N177);
nor NOR4 (N1084, N1080, N1042, N390, N116);
or OR2 (N1085, N1073, N960);
and AND4 (N1086, N1081, N712, N910, N137);
buf BUF1 (N1087, N1083);
nor NOR4 (N1088, N1057, N741, N403, N663);
nand NAND4 (N1089, N1082, N1034, N155, N599);
xor XOR2 (N1090, N1085, N1055);
xor XOR2 (N1091, N1072, N410);
not NOT1 (N1092, N1070);
xor XOR2 (N1093, N1086, N62);
and AND3 (N1094, N1087, N705, N582);
not NOT1 (N1095, N1078);
and AND3 (N1096, N1089, N916, N215);
xor XOR2 (N1097, N1075, N909);
and AND2 (N1098, N1094, N490);
not NOT1 (N1099, N1096);
or OR4 (N1100, N1099, N917, N360, N652);
not NOT1 (N1101, N1088);
buf BUF1 (N1102, N1091);
buf BUF1 (N1103, N1092);
and AND4 (N1104, N1084, N478, N1064, N181);
and AND3 (N1105, N1101, N595, N1015);
nor NOR3 (N1106, N1105, N1054, N494);
xor XOR2 (N1107, N1090, N172);
xor XOR2 (N1108, N1097, N511);
not NOT1 (N1109, N1100);
or OR3 (N1110, N1109, N602, N599);
and AND3 (N1111, N1110, N306, N273);
not NOT1 (N1112, N1102);
nand NAND2 (N1113, N1108, N909);
buf BUF1 (N1114, N1106);
not NOT1 (N1115, N1093);
buf BUF1 (N1116, N1107);
and AND3 (N1117, N1115, N407, N327);
xor XOR2 (N1118, N1114, N70);
buf BUF1 (N1119, N1113);
xor XOR2 (N1120, N1112, N614);
nor NOR4 (N1121, N1095, N876, N128, N1037);
or OR2 (N1122, N1119, N105);
not NOT1 (N1123, N1103);
or OR3 (N1124, N1118, N400, N325);
buf BUF1 (N1125, N1111);
nand NAND3 (N1126, N1124, N579, N310);
nand NAND2 (N1127, N1121, N172);
not NOT1 (N1128, N1117);
not NOT1 (N1129, N1125);
xor XOR2 (N1130, N1122, N967);
or OR4 (N1131, N1126, N118, N873, N1023);
and AND2 (N1132, N1104, N561);
buf BUF1 (N1133, N1127);
nor NOR3 (N1134, N1123, N977, N94);
nor NOR3 (N1135, N1128, N721, N554);
not NOT1 (N1136, N1130);
not NOT1 (N1137, N1131);
or OR2 (N1138, N1120, N495);
buf BUF1 (N1139, N1133);
and AND2 (N1140, N1137, N197);
nand NAND2 (N1141, N1129, N52);
nor NOR2 (N1142, N1136, N377);
buf BUF1 (N1143, N1132);
xor XOR2 (N1144, N1138, N890);
or OR3 (N1145, N1142, N506, N786);
nand NAND3 (N1146, N1141, N70, N609);
and AND4 (N1147, N1146, N1065, N791, N341);
not NOT1 (N1148, N1143);
buf BUF1 (N1149, N1139);
nor NOR2 (N1150, N1144, N1131);
buf BUF1 (N1151, N1140);
buf BUF1 (N1152, N1149);
xor XOR2 (N1153, N1152, N294);
or OR2 (N1154, N1151, N296);
nand NAND4 (N1155, N1147, N710, N726, N909);
nand NAND4 (N1156, N1153, N1111, N928, N372);
or OR4 (N1157, N1134, N348, N118, N230);
xor XOR2 (N1158, N1116, N232);
nor NOR4 (N1159, N1135, N1082, N488, N493);
or OR2 (N1160, N1156, N1093);
or OR4 (N1161, N1145, N204, N556, N356);
nor NOR3 (N1162, N1157, N96, N920);
or OR3 (N1163, N1161, N797, N112);
nand NAND4 (N1164, N1158, N1156, N151, N877);
nand NAND2 (N1165, N1148, N1032);
xor XOR2 (N1166, N1163, N1116);
nor NOR4 (N1167, N1160, N740, N962, N286);
xor XOR2 (N1168, N1154, N625);
not NOT1 (N1169, N1098);
nor NOR3 (N1170, N1164, N240, N197);
not NOT1 (N1171, N1162);
or OR3 (N1172, N1165, N305, N853);
nor NOR4 (N1173, N1168, N1022, N306, N46);
buf BUF1 (N1174, N1173);
nand NAND2 (N1175, N1169, N869);
or OR3 (N1176, N1155, N1159, N277);
xor XOR2 (N1177, N268, N955);
xor XOR2 (N1178, N1176, N443);
nor NOR2 (N1179, N1150, N873);
xor XOR2 (N1180, N1174, N372);
nor NOR2 (N1181, N1180, N874);
nor NOR2 (N1182, N1178, N1053);
or OR2 (N1183, N1170, N133);
nor NOR3 (N1184, N1167, N606, N271);
not NOT1 (N1185, N1172);
not NOT1 (N1186, N1175);
not NOT1 (N1187, N1183);
buf BUF1 (N1188, N1171);
and AND3 (N1189, N1177, N916, N237);
buf BUF1 (N1190, N1179);
xor XOR2 (N1191, N1184, N985);
xor XOR2 (N1192, N1185, N908);
xor XOR2 (N1193, N1182, N263);
xor XOR2 (N1194, N1166, N170);
nor NOR4 (N1195, N1193, N1065, N1176, N930);
nand NAND2 (N1196, N1190, N35);
and AND2 (N1197, N1195, N1136);
xor XOR2 (N1198, N1196, N440);
nor NOR2 (N1199, N1186, N1055);
or OR2 (N1200, N1187, N999);
or OR3 (N1201, N1188, N207, N1157);
buf BUF1 (N1202, N1181);
xor XOR2 (N1203, N1201, N140);
not NOT1 (N1204, N1203);
buf BUF1 (N1205, N1198);
and AND4 (N1206, N1194, N502, N243, N12);
xor XOR2 (N1207, N1199, N65);
buf BUF1 (N1208, N1192);
not NOT1 (N1209, N1205);
buf BUF1 (N1210, N1202);
or OR3 (N1211, N1207, N18, N426);
and AND3 (N1212, N1206, N514, N889);
nand NAND2 (N1213, N1197, N66);
nand NAND2 (N1214, N1212, N1049);
not NOT1 (N1215, N1204);
xor XOR2 (N1216, N1210, N348);
or OR2 (N1217, N1215, N1018);
buf BUF1 (N1218, N1191);
or OR4 (N1219, N1214, N241, N936, N539);
not NOT1 (N1220, N1208);
xor XOR2 (N1221, N1218, N579);
or OR2 (N1222, N1209, N429);
not NOT1 (N1223, N1211);
nand NAND3 (N1224, N1216, N85, N588);
nor NOR2 (N1225, N1224, N888);
xor XOR2 (N1226, N1220, N308);
xor XOR2 (N1227, N1222, N213);
buf BUF1 (N1228, N1223);
nor NOR2 (N1229, N1213, N292);
or OR3 (N1230, N1219, N110, N467);
nand NAND3 (N1231, N1230, N229, N1161);
nor NOR2 (N1232, N1225, N176);
xor XOR2 (N1233, N1229, N646);
or OR2 (N1234, N1189, N891);
nand NAND2 (N1235, N1233, N1185);
not NOT1 (N1236, N1227);
buf BUF1 (N1237, N1232);
buf BUF1 (N1238, N1237);
buf BUF1 (N1239, N1236);
and AND4 (N1240, N1228, N974, N125, N72);
nor NOR2 (N1241, N1231, N857);
buf BUF1 (N1242, N1200);
and AND2 (N1243, N1239, N690);
or OR4 (N1244, N1240, N140, N140, N960);
and AND3 (N1245, N1221, N979, N489);
nor NOR3 (N1246, N1234, N102, N1131);
and AND3 (N1247, N1241, N670, N597);
nand NAND3 (N1248, N1217, N567, N415);
and AND3 (N1249, N1244, N475, N837);
nor NOR2 (N1250, N1246, N1);
nor NOR3 (N1251, N1248, N1154, N809);
not NOT1 (N1252, N1249);
nand NAND4 (N1253, N1235, N627, N595, N49);
xor XOR2 (N1254, N1245, N112);
or OR2 (N1255, N1250, N783);
buf BUF1 (N1256, N1255);
nand NAND4 (N1257, N1247, N1242, N274, N295);
or OR4 (N1258, N413, N11, N474, N612);
or OR3 (N1259, N1252, N1005, N742);
nor NOR2 (N1260, N1254, N37);
nand NAND2 (N1261, N1256, N1099);
or OR2 (N1262, N1260, N326);
xor XOR2 (N1263, N1253, N704);
and AND2 (N1264, N1258, N65);
nor NOR2 (N1265, N1226, N108);
xor XOR2 (N1266, N1243, N1157);
or OR4 (N1267, N1259, N566, N193, N826);
or OR3 (N1268, N1263, N1199, N517);
or OR3 (N1269, N1264, N1199, N840);
buf BUF1 (N1270, N1267);
buf BUF1 (N1271, N1270);
and AND3 (N1272, N1271, N399, N592);
xor XOR2 (N1273, N1269, N737);
and AND4 (N1274, N1266, N1123, N1096, N25);
not NOT1 (N1275, N1261);
buf BUF1 (N1276, N1238);
not NOT1 (N1277, N1262);
xor XOR2 (N1278, N1274, N761);
nor NOR2 (N1279, N1277, N39);
nand NAND4 (N1280, N1275, N1122, N271, N1101);
and AND3 (N1281, N1251, N467, N699);
nor NOR4 (N1282, N1272, N284, N220, N994);
buf BUF1 (N1283, N1280);
nor NOR2 (N1284, N1268, N1260);
nand NAND3 (N1285, N1276, N1182, N254);
nand NAND2 (N1286, N1265, N452);
buf BUF1 (N1287, N1283);
nor NOR3 (N1288, N1287, N651, N53);
xor XOR2 (N1289, N1282, N851);
not NOT1 (N1290, N1289);
nand NAND3 (N1291, N1285, N311, N484);
nor NOR3 (N1292, N1257, N62, N88);
nor NOR2 (N1293, N1278, N602);
not NOT1 (N1294, N1273);
buf BUF1 (N1295, N1291);
nor NOR3 (N1296, N1292, N359, N374);
not NOT1 (N1297, N1286);
buf BUF1 (N1298, N1279);
buf BUF1 (N1299, N1298);
buf BUF1 (N1300, N1288);
xor XOR2 (N1301, N1299, N275);
or OR3 (N1302, N1281, N66, N356);
buf BUF1 (N1303, N1284);
xor XOR2 (N1304, N1301, N11);
nor NOR3 (N1305, N1296, N417, N1149);
or OR3 (N1306, N1294, N982, N843);
nand NAND3 (N1307, N1300, N347, N73);
buf BUF1 (N1308, N1295);
buf BUF1 (N1309, N1293);
or OR2 (N1310, N1297, N904);
nand NAND4 (N1311, N1290, N851, N567, N1030);
nor NOR4 (N1312, N1311, N1140, N431, N677);
and AND4 (N1313, N1309, N1025, N700, N720);
and AND3 (N1314, N1302, N487, N857);
xor XOR2 (N1315, N1304, N372);
xor XOR2 (N1316, N1313, N754);
not NOT1 (N1317, N1303);
nor NOR2 (N1318, N1305, N307);
not NOT1 (N1319, N1315);
or OR4 (N1320, N1318, N1262, N1022, N381);
and AND3 (N1321, N1320, N857, N723);
and AND3 (N1322, N1310, N678, N843);
not NOT1 (N1323, N1321);
and AND3 (N1324, N1314, N533, N135);
buf BUF1 (N1325, N1319);
and AND2 (N1326, N1317, N781);
buf BUF1 (N1327, N1322);
not NOT1 (N1328, N1308);
and AND3 (N1329, N1307, N122, N389);
or OR4 (N1330, N1326, N284, N615, N913);
or OR4 (N1331, N1325, N1075, N89, N316);
buf BUF1 (N1332, N1323);
or OR3 (N1333, N1316, N193, N492);
xor XOR2 (N1334, N1331, N1066);
not NOT1 (N1335, N1328);
nand NAND2 (N1336, N1329, N944);
not NOT1 (N1337, N1324);
xor XOR2 (N1338, N1336, N595);
nand NAND4 (N1339, N1333, N1177, N453, N1292);
buf BUF1 (N1340, N1339);
or OR4 (N1341, N1332, N106, N49, N388);
buf BUF1 (N1342, N1334);
or OR2 (N1343, N1306, N691);
nor NOR2 (N1344, N1338, N185);
nand NAND4 (N1345, N1335, N131, N401, N1071);
or OR2 (N1346, N1343, N981);
or OR3 (N1347, N1312, N905, N1069);
and AND2 (N1348, N1327, N436);
nor NOR3 (N1349, N1337, N71, N495);
and AND2 (N1350, N1347, N596);
xor XOR2 (N1351, N1345, N751);
buf BUF1 (N1352, N1342);
or OR4 (N1353, N1341, N1024, N945, N791);
or OR2 (N1354, N1346, N502);
not NOT1 (N1355, N1348);
nand NAND4 (N1356, N1352, N893, N66, N300);
xor XOR2 (N1357, N1330, N6);
xor XOR2 (N1358, N1344, N322);
xor XOR2 (N1359, N1357, N445);
or OR4 (N1360, N1359, N108, N1265, N1059);
nand NAND4 (N1361, N1349, N225, N438, N1138);
and AND4 (N1362, N1360, N622, N1223, N33);
or OR2 (N1363, N1353, N699);
nand NAND4 (N1364, N1355, N1022, N689, N869);
nand NAND3 (N1365, N1351, N425, N216);
buf BUF1 (N1366, N1365);
nand NAND4 (N1367, N1358, N290, N452, N691);
or OR2 (N1368, N1350, N1223);
xor XOR2 (N1369, N1367, N441);
or OR4 (N1370, N1354, N226, N1197, N1261);
xor XOR2 (N1371, N1340, N521);
not NOT1 (N1372, N1363);
and AND3 (N1373, N1362, N1009, N952);
xor XOR2 (N1374, N1368, N243);
xor XOR2 (N1375, N1366, N287);
or OR4 (N1376, N1373, N800, N144, N1244);
and AND4 (N1377, N1370, N1207, N798, N1139);
not NOT1 (N1378, N1376);
xor XOR2 (N1379, N1377, N675);
nand NAND3 (N1380, N1379, N109, N828);
not NOT1 (N1381, N1380);
buf BUF1 (N1382, N1374);
or OR4 (N1383, N1378, N343, N644, N759);
buf BUF1 (N1384, N1383);
xor XOR2 (N1385, N1384, N1230);
nor NOR3 (N1386, N1364, N799, N496);
buf BUF1 (N1387, N1361);
and AND4 (N1388, N1356, N804, N271, N210);
and AND3 (N1389, N1387, N193, N129);
not NOT1 (N1390, N1385);
buf BUF1 (N1391, N1372);
not NOT1 (N1392, N1371);
or OR2 (N1393, N1389, N1205);
or OR4 (N1394, N1369, N880, N94, N671);
or OR4 (N1395, N1382, N740, N590, N324);
not NOT1 (N1396, N1388);
not NOT1 (N1397, N1375);
nor NOR2 (N1398, N1397, N103);
nor NOR3 (N1399, N1398, N957, N887);
xor XOR2 (N1400, N1392, N1165);
nor NOR2 (N1401, N1395, N1395);
nor NOR3 (N1402, N1390, N597, N1031);
nor NOR3 (N1403, N1400, N667, N550);
or OR2 (N1404, N1402, N809);
nand NAND4 (N1405, N1396, N150, N1036, N1367);
or OR2 (N1406, N1393, N1323);
not NOT1 (N1407, N1404);
or OR2 (N1408, N1401, N879);
not NOT1 (N1409, N1381);
not NOT1 (N1410, N1409);
or OR2 (N1411, N1407, N681);
and AND2 (N1412, N1399, N458);
nand NAND3 (N1413, N1410, N1049, N1228);
and AND4 (N1414, N1413, N325, N1243, N985);
and AND3 (N1415, N1394, N1126, N240);
and AND2 (N1416, N1411, N876);
or OR4 (N1417, N1414, N770, N61, N1161);
buf BUF1 (N1418, N1417);
not NOT1 (N1419, N1403);
nand NAND3 (N1420, N1406, N1087, N904);
not NOT1 (N1421, N1420);
buf BUF1 (N1422, N1412);
nand NAND3 (N1423, N1386, N497, N612);
nand NAND3 (N1424, N1391, N642, N954);
or OR3 (N1425, N1424, N789, N313);
nor NOR4 (N1426, N1408, N1000, N1222, N206);
nor NOR3 (N1427, N1415, N1015, N1026);
and AND4 (N1428, N1419, N1151, N499, N1192);
and AND3 (N1429, N1427, N162, N1173);
and AND4 (N1430, N1428, N51, N1105, N331);
xor XOR2 (N1431, N1429, N70);
not NOT1 (N1432, N1405);
or OR2 (N1433, N1416, N1374);
buf BUF1 (N1434, N1422);
buf BUF1 (N1435, N1418);
nand NAND3 (N1436, N1433, N416, N508);
and AND2 (N1437, N1423, N991);
and AND2 (N1438, N1431, N1373);
or OR2 (N1439, N1426, N1384);
and AND3 (N1440, N1425, N142, N1396);
buf BUF1 (N1441, N1435);
nand NAND3 (N1442, N1432, N461, N423);
nor NOR4 (N1443, N1439, N761, N561, N1239);
buf BUF1 (N1444, N1443);
not NOT1 (N1445, N1442);
nor NOR3 (N1446, N1437, N1159, N213);
and AND3 (N1447, N1421, N757, N252);
and AND2 (N1448, N1430, N255);
buf BUF1 (N1449, N1448);
and AND4 (N1450, N1445, N1354, N1204, N223);
nand NAND4 (N1451, N1438, N383, N159, N1361);
xor XOR2 (N1452, N1436, N461);
buf BUF1 (N1453, N1440);
not NOT1 (N1454, N1447);
xor XOR2 (N1455, N1446, N49);
nor NOR2 (N1456, N1444, N1429);
xor XOR2 (N1457, N1453, N375);
xor XOR2 (N1458, N1452, N411);
xor XOR2 (N1459, N1449, N757);
and AND4 (N1460, N1434, N1011, N699, N587);
buf BUF1 (N1461, N1455);
nor NOR3 (N1462, N1460, N151, N372);
buf BUF1 (N1463, N1461);
or OR3 (N1464, N1451, N357, N690);
nand NAND2 (N1465, N1450, N834);
and AND2 (N1466, N1457, N1249);
nand NAND4 (N1467, N1464, N1384, N36, N426);
not NOT1 (N1468, N1465);
and AND3 (N1469, N1458, N1229, N1168);
buf BUF1 (N1470, N1469);
or OR4 (N1471, N1459, N812, N985, N64);
nand NAND4 (N1472, N1441, N510, N1054, N402);
or OR4 (N1473, N1454, N249, N379, N185);
or OR2 (N1474, N1473, N179);
buf BUF1 (N1475, N1467);
nor NOR4 (N1476, N1466, N690, N463, N1428);
nor NOR2 (N1477, N1471, N968);
and AND4 (N1478, N1476, N897, N246, N1455);
not NOT1 (N1479, N1456);
or OR4 (N1480, N1479, N806, N746, N1373);
not NOT1 (N1481, N1478);
not NOT1 (N1482, N1480);
xor XOR2 (N1483, N1463, N1298);
nand NAND2 (N1484, N1474, N537);
or OR4 (N1485, N1482, N366, N132, N809);
nand NAND4 (N1486, N1477, N713, N1280, N1000);
and AND3 (N1487, N1481, N228, N386);
xor XOR2 (N1488, N1468, N595);
not NOT1 (N1489, N1484);
or OR3 (N1490, N1487, N116, N981);
not NOT1 (N1491, N1470);
not NOT1 (N1492, N1485);
not NOT1 (N1493, N1462);
or OR4 (N1494, N1489, N1080, N1065, N1471);
buf BUF1 (N1495, N1493);
or OR2 (N1496, N1491, N1278);
or OR3 (N1497, N1475, N1127, N34);
nor NOR3 (N1498, N1488, N749, N47);
or OR2 (N1499, N1486, N1169);
and AND3 (N1500, N1497, N268, N186);
xor XOR2 (N1501, N1483, N1039);
xor XOR2 (N1502, N1498, N1084);
xor XOR2 (N1503, N1496, N660);
and AND2 (N1504, N1499, N546);
buf BUF1 (N1505, N1504);
nand NAND2 (N1506, N1490, N1443);
nand NAND3 (N1507, N1495, N998, N704);
and AND3 (N1508, N1472, N1348, N1132);
not NOT1 (N1509, N1503);
nor NOR2 (N1510, N1507, N1010);
or OR2 (N1511, N1510, N1358);
nor NOR2 (N1512, N1500, N196);
not NOT1 (N1513, N1506);
buf BUF1 (N1514, N1492);
nand NAND4 (N1515, N1514, N430, N542, N1039);
not NOT1 (N1516, N1502);
nor NOR2 (N1517, N1516, N517);
nor NOR2 (N1518, N1505, N128);
nand NAND2 (N1519, N1494, N1408);
nand NAND4 (N1520, N1501, N89, N533, N669);
or OR3 (N1521, N1515, N20, N983);
and AND4 (N1522, N1521, N925, N686, N803);
not NOT1 (N1523, N1513);
buf BUF1 (N1524, N1518);
nor NOR4 (N1525, N1508, N9, N1049, N20);
and AND3 (N1526, N1509, N1426, N1447);
nand NAND2 (N1527, N1524, N128);
or OR4 (N1528, N1512, N326, N1274, N1198);
xor XOR2 (N1529, N1526, N584);
or OR4 (N1530, N1523, N1492, N838, N822);
or OR2 (N1531, N1520, N1420);
or OR4 (N1532, N1522, N1266, N734, N1357);
and AND4 (N1533, N1511, N625, N1023, N1515);
or OR3 (N1534, N1531, N723, N380);
not NOT1 (N1535, N1532);
not NOT1 (N1536, N1519);
buf BUF1 (N1537, N1529);
buf BUF1 (N1538, N1534);
xor XOR2 (N1539, N1517, N742);
or OR4 (N1540, N1528, N454, N561, N499);
not NOT1 (N1541, N1535);
not NOT1 (N1542, N1527);
and AND3 (N1543, N1537, N48, N1496);
nor NOR3 (N1544, N1539, N597, N153);
not NOT1 (N1545, N1538);
nand NAND2 (N1546, N1545, N346);
not NOT1 (N1547, N1536);
or OR4 (N1548, N1533, N564, N750, N81);
nand NAND3 (N1549, N1542, N1098, N435);
not NOT1 (N1550, N1530);
or OR3 (N1551, N1543, N614, N1323);
not NOT1 (N1552, N1550);
nand NAND2 (N1553, N1540, N1152);
xor XOR2 (N1554, N1541, N698);
nand NAND2 (N1555, N1547, N1301);
nor NOR2 (N1556, N1554, N194);
xor XOR2 (N1557, N1544, N1153);
not NOT1 (N1558, N1553);
xor XOR2 (N1559, N1546, N1260);
xor XOR2 (N1560, N1549, N308);
and AND3 (N1561, N1556, N358, N380);
and AND4 (N1562, N1560, N154, N1075, N1514);
buf BUF1 (N1563, N1561);
and AND4 (N1564, N1557, N679, N1077, N470);
or OR2 (N1565, N1559, N251);
xor XOR2 (N1566, N1551, N1106);
xor XOR2 (N1567, N1525, N410);
and AND4 (N1568, N1548, N1253, N1237, N620);
or OR3 (N1569, N1566, N1057, N1137);
or OR4 (N1570, N1567, N1444, N902, N802);
and AND4 (N1571, N1563, N693, N186, N468);
buf BUF1 (N1572, N1569);
and AND4 (N1573, N1570, N701, N188, N850);
nor NOR4 (N1574, N1564, N83, N1530, N255);
or OR2 (N1575, N1562, N922);
xor XOR2 (N1576, N1558, N632);
or OR3 (N1577, N1575, N1337, N220);
and AND3 (N1578, N1568, N385, N704);
or OR4 (N1579, N1565, N1541, N253, N186);
nand NAND4 (N1580, N1574, N538, N603, N208);
buf BUF1 (N1581, N1580);
nor NOR3 (N1582, N1577, N1035, N1562);
nor NOR2 (N1583, N1576, N1096);
or OR2 (N1584, N1578, N727);
not NOT1 (N1585, N1552);
or OR4 (N1586, N1581, N682, N1152, N1110);
nand NAND2 (N1587, N1572, N363);
nand NAND2 (N1588, N1582, N251);
or OR3 (N1589, N1585, N541, N726);
or OR4 (N1590, N1586, N1450, N815, N316);
nor NOR3 (N1591, N1555, N1318, N204);
nand NAND4 (N1592, N1579, N276, N1075, N69);
nor NOR4 (N1593, N1591, N435, N1543, N1520);
not NOT1 (N1594, N1573);
nand NAND2 (N1595, N1593, N853);
nand NAND3 (N1596, N1594, N88, N1550);
or OR2 (N1597, N1587, N1109);
not NOT1 (N1598, N1592);
nand NAND2 (N1599, N1590, N954);
not NOT1 (N1600, N1571);
not NOT1 (N1601, N1588);
nor NOR3 (N1602, N1596, N1042, N1582);
nor NOR3 (N1603, N1583, N1586, N202);
or OR3 (N1604, N1597, N611, N348);
nand NAND3 (N1605, N1598, N343, N1308);
buf BUF1 (N1606, N1600);
and AND4 (N1607, N1595, N64, N1482, N373);
xor XOR2 (N1608, N1589, N687);
or OR4 (N1609, N1599, N1327, N60, N507);
or OR2 (N1610, N1584, N336);
nand NAND3 (N1611, N1603, N790, N1046);
not NOT1 (N1612, N1601);
nor NOR4 (N1613, N1612, N584, N1303, N760);
nand NAND3 (N1614, N1605, N1186, N943);
nor NOR3 (N1615, N1609, N280, N429);
xor XOR2 (N1616, N1608, N1343);
buf BUF1 (N1617, N1610);
nor NOR3 (N1618, N1617, N1223, N1471);
or OR3 (N1619, N1602, N29, N1467);
not NOT1 (N1620, N1619);
xor XOR2 (N1621, N1607, N973);
nand NAND3 (N1622, N1621, N948, N539);
buf BUF1 (N1623, N1611);
and AND4 (N1624, N1620, N358, N67, N412);
buf BUF1 (N1625, N1613);
and AND4 (N1626, N1616, N1035, N982, N833);
buf BUF1 (N1627, N1604);
buf BUF1 (N1628, N1625);
not NOT1 (N1629, N1626);
buf BUF1 (N1630, N1606);
xor XOR2 (N1631, N1622, N1035);
and AND2 (N1632, N1623, N988);
and AND3 (N1633, N1631, N828, N885);
xor XOR2 (N1634, N1614, N504);
and AND4 (N1635, N1634, N936, N1131, N101);
nor NOR3 (N1636, N1629, N789, N78);
nand NAND4 (N1637, N1615, N1043, N257, N174);
xor XOR2 (N1638, N1628, N503);
nand NAND2 (N1639, N1635, N1106);
not NOT1 (N1640, N1624);
or OR4 (N1641, N1636, N3, N1375, N523);
not NOT1 (N1642, N1640);
or OR4 (N1643, N1637, N622, N331, N500);
not NOT1 (N1644, N1643);
nand NAND2 (N1645, N1633, N1465);
and AND4 (N1646, N1638, N1301, N1, N211);
and AND4 (N1647, N1642, N281, N326, N1276);
buf BUF1 (N1648, N1647);
xor XOR2 (N1649, N1646, N1132);
not NOT1 (N1650, N1649);
buf BUF1 (N1651, N1648);
buf BUF1 (N1652, N1641);
xor XOR2 (N1653, N1630, N807);
nor NOR2 (N1654, N1653, N425);
nand NAND2 (N1655, N1651, N141);
xor XOR2 (N1656, N1654, N561);
or OR2 (N1657, N1656, N1483);
not NOT1 (N1658, N1655);
nor NOR4 (N1659, N1650, N1171, N409, N24);
nor NOR2 (N1660, N1627, N10);
buf BUF1 (N1661, N1660);
or OR2 (N1662, N1618, N1156);
xor XOR2 (N1663, N1662, N1127);
nor NOR3 (N1664, N1639, N176, N135);
and AND3 (N1665, N1644, N967, N513);
nor NOR2 (N1666, N1664, N378);
nand NAND2 (N1667, N1657, N787);
xor XOR2 (N1668, N1665, N817);
buf BUF1 (N1669, N1668);
buf BUF1 (N1670, N1667);
xor XOR2 (N1671, N1661, N22);
nand NAND2 (N1672, N1670, N725);
and AND2 (N1673, N1671, N340);
not NOT1 (N1674, N1659);
or OR3 (N1675, N1673, N129, N1381);
buf BUF1 (N1676, N1652);
and AND4 (N1677, N1658, N700, N1487, N372);
buf BUF1 (N1678, N1669);
nand NAND3 (N1679, N1663, N189, N959);
not NOT1 (N1680, N1677);
and AND4 (N1681, N1666, N734, N1278, N494);
nand NAND2 (N1682, N1678, N767);
buf BUF1 (N1683, N1674);
or OR3 (N1684, N1672, N1437, N1017);
not NOT1 (N1685, N1684);
and AND4 (N1686, N1676, N1578, N207, N887);
not NOT1 (N1687, N1675);
buf BUF1 (N1688, N1681);
not NOT1 (N1689, N1687);
nor NOR3 (N1690, N1683, N448, N374);
buf BUF1 (N1691, N1686);
and AND3 (N1692, N1691, N425, N1379);
buf BUF1 (N1693, N1680);
nor NOR3 (N1694, N1679, N1334, N636);
nand NAND3 (N1695, N1689, N159, N1033);
and AND2 (N1696, N1693, N126);
nor NOR2 (N1697, N1632, N828);
not NOT1 (N1698, N1696);
xor XOR2 (N1699, N1695, N623);
not NOT1 (N1700, N1682);
or OR4 (N1701, N1690, N980, N1160, N1320);
and AND2 (N1702, N1694, N1288);
or OR3 (N1703, N1645, N256, N206);
buf BUF1 (N1704, N1699);
xor XOR2 (N1705, N1702, N1348);
buf BUF1 (N1706, N1698);
xor XOR2 (N1707, N1697, N1691);
nand NAND3 (N1708, N1685, N644, N1262);
nand NAND2 (N1709, N1708, N30);
xor XOR2 (N1710, N1706, N641);
nor NOR3 (N1711, N1704, N844, N368);
and AND4 (N1712, N1709, N1318, N965, N14);
not NOT1 (N1713, N1707);
not NOT1 (N1714, N1688);
nand NAND3 (N1715, N1705, N71, N790);
not NOT1 (N1716, N1701);
nor NOR3 (N1717, N1714, N227, N1197);
buf BUF1 (N1718, N1703);
buf BUF1 (N1719, N1716);
buf BUF1 (N1720, N1717);
not NOT1 (N1721, N1720);
buf BUF1 (N1722, N1713);
nor NOR2 (N1723, N1721, N1490);
or OR3 (N1724, N1722, N457, N1306);
xor XOR2 (N1725, N1692, N818);
buf BUF1 (N1726, N1719);
buf BUF1 (N1727, N1725);
not NOT1 (N1728, N1727);
nand NAND3 (N1729, N1700, N179, N246);
xor XOR2 (N1730, N1712, N605);
buf BUF1 (N1731, N1710);
nor NOR2 (N1732, N1715, N1488);
xor XOR2 (N1733, N1731, N860);
buf BUF1 (N1734, N1733);
nor NOR2 (N1735, N1730, N207);
nand NAND4 (N1736, N1723, N1725, N1548, N913);
or OR2 (N1737, N1711, N619);
buf BUF1 (N1738, N1728);
and AND3 (N1739, N1738, N1173, N1464);
not NOT1 (N1740, N1737);
nor NOR3 (N1741, N1734, N772, N227);
nand NAND2 (N1742, N1718, N1618);
xor XOR2 (N1743, N1735, N346);
buf BUF1 (N1744, N1742);
nand NAND4 (N1745, N1743, N1521, N1502, N1442);
nor NOR2 (N1746, N1744, N838);
and AND4 (N1747, N1729, N1453, N800, N1411);
nand NAND4 (N1748, N1747, N439, N358, N1580);
not NOT1 (N1749, N1745);
nor NOR4 (N1750, N1726, N1247, N1402, N909);
buf BUF1 (N1751, N1732);
or OR4 (N1752, N1739, N972, N1695, N785);
nand NAND2 (N1753, N1724, N1220);
and AND4 (N1754, N1753, N1208, N1586, N1274);
not NOT1 (N1755, N1752);
buf BUF1 (N1756, N1746);
xor XOR2 (N1757, N1754, N1658);
or OR4 (N1758, N1757, N1700, N161, N19);
or OR2 (N1759, N1750, N529);
xor XOR2 (N1760, N1755, N1460);
nor NOR4 (N1761, N1740, N434, N675, N402);
and AND3 (N1762, N1736, N1515, N251);
xor XOR2 (N1763, N1759, N1330);
xor XOR2 (N1764, N1762, N646);
and AND4 (N1765, N1748, N655, N1726, N1230);
not NOT1 (N1766, N1761);
and AND4 (N1767, N1758, N846, N1532, N997);
or OR2 (N1768, N1749, N349);
and AND2 (N1769, N1766, N449);
xor XOR2 (N1770, N1768, N304);
and AND4 (N1771, N1767, N904, N958, N1337);
and AND2 (N1772, N1760, N33);
xor XOR2 (N1773, N1751, N1618);
xor XOR2 (N1774, N1770, N523);
xor XOR2 (N1775, N1774, N157);
nand NAND4 (N1776, N1741, N997, N1691, N1396);
nor NOR4 (N1777, N1756, N121, N85, N208);
not NOT1 (N1778, N1772);
nor NOR2 (N1779, N1777, N566);
or OR2 (N1780, N1764, N510);
not NOT1 (N1781, N1778);
not NOT1 (N1782, N1776);
xor XOR2 (N1783, N1779, N1476);
and AND2 (N1784, N1781, N260);
xor XOR2 (N1785, N1769, N5);
xor XOR2 (N1786, N1784, N1288);
or OR4 (N1787, N1771, N889, N332, N972);
nand NAND4 (N1788, N1787, N502, N951, N253);
and AND2 (N1789, N1780, N1227);
xor XOR2 (N1790, N1785, N198);
or OR2 (N1791, N1775, N673);
or OR4 (N1792, N1789, N1585, N587, N1614);
nor NOR2 (N1793, N1786, N1139);
or OR4 (N1794, N1793, N1098, N137, N431);
nand NAND3 (N1795, N1794, N385, N639);
buf BUF1 (N1796, N1765);
nand NAND2 (N1797, N1763, N431);
xor XOR2 (N1798, N1797, N325);
nor NOR2 (N1799, N1796, N1336);
not NOT1 (N1800, N1795);
or OR4 (N1801, N1782, N1623, N1036, N92);
buf BUF1 (N1802, N1801);
nand NAND2 (N1803, N1773, N1774);
or OR3 (N1804, N1788, N1064, N1766);
buf BUF1 (N1805, N1791);
nor NOR4 (N1806, N1802, N1555, N904, N996);
and AND4 (N1807, N1800, N100, N962, N240);
not NOT1 (N1808, N1783);
nand NAND3 (N1809, N1804, N444, N206);
or OR2 (N1810, N1809, N985);
buf BUF1 (N1811, N1790);
or OR4 (N1812, N1810, N199, N660, N188);
buf BUF1 (N1813, N1803);
nand NAND2 (N1814, N1792, N1153);
nor NOR3 (N1815, N1813, N1131, N1601);
nor NOR3 (N1816, N1807, N105, N1385);
or OR3 (N1817, N1805, N220, N310);
not NOT1 (N1818, N1816);
nand NAND3 (N1819, N1799, N264, N808);
nand NAND2 (N1820, N1818, N1563);
not NOT1 (N1821, N1812);
buf BUF1 (N1822, N1819);
nand NAND2 (N1823, N1822, N1329);
nand NAND4 (N1824, N1806, N1161, N681, N1106);
not NOT1 (N1825, N1814);
and AND3 (N1826, N1824, N87, N855);
not NOT1 (N1827, N1811);
xor XOR2 (N1828, N1817, N1605);
or OR4 (N1829, N1820, N301, N849, N18);
not NOT1 (N1830, N1829);
or OR3 (N1831, N1821, N51, N1093);
or OR2 (N1832, N1827, N1705);
not NOT1 (N1833, N1823);
not NOT1 (N1834, N1826);
xor XOR2 (N1835, N1834, N1436);
and AND4 (N1836, N1832, N1463, N1072, N1089);
or OR2 (N1837, N1836, N1135);
nand NAND3 (N1838, N1798, N378, N610);
buf BUF1 (N1839, N1815);
not NOT1 (N1840, N1828);
nand NAND3 (N1841, N1833, N48, N1476);
not NOT1 (N1842, N1839);
or OR3 (N1843, N1831, N749, N1494);
nand NAND4 (N1844, N1837, N233, N1283, N1441);
xor XOR2 (N1845, N1835, N783);
buf BUF1 (N1846, N1841);
nor NOR3 (N1847, N1846, N46, N207);
and AND2 (N1848, N1808, N1107);
nor NOR2 (N1849, N1842, N468);
and AND3 (N1850, N1838, N284, N402);
and AND4 (N1851, N1843, N29, N636, N522);
xor XOR2 (N1852, N1851, N441);
nand NAND3 (N1853, N1844, N390, N1345);
nand NAND4 (N1854, N1852, N645, N722, N157);
nor NOR2 (N1855, N1849, N832);
nand NAND3 (N1856, N1855, N332, N1819);
nor NOR4 (N1857, N1856, N355, N1799, N149);
not NOT1 (N1858, N1845);
not NOT1 (N1859, N1850);
nand NAND4 (N1860, N1825, N842, N598, N953);
buf BUF1 (N1861, N1859);
and AND2 (N1862, N1830, N212);
buf BUF1 (N1863, N1862);
buf BUF1 (N1864, N1861);
nand NAND3 (N1865, N1847, N895, N22);
nor NOR4 (N1866, N1840, N975, N624, N532);
nor NOR3 (N1867, N1860, N297, N474);
buf BUF1 (N1868, N1867);
and AND3 (N1869, N1853, N502, N923);
or OR4 (N1870, N1858, N1258, N1515, N86);
nor NOR4 (N1871, N1848, N746, N330, N958);
or OR2 (N1872, N1868, N1441);
xor XOR2 (N1873, N1857, N903);
xor XOR2 (N1874, N1872, N585);
xor XOR2 (N1875, N1874, N851);
xor XOR2 (N1876, N1863, N651);
nor NOR4 (N1877, N1870, N1557, N576, N81);
nand NAND3 (N1878, N1865, N193, N492);
xor XOR2 (N1879, N1877, N1794);
and AND4 (N1880, N1866, N1687, N14, N1514);
xor XOR2 (N1881, N1875, N1625);
nor NOR3 (N1882, N1878, N456, N1772);
or OR2 (N1883, N1869, N283);
or OR2 (N1884, N1864, N1680);
xor XOR2 (N1885, N1880, N448);
nand NAND4 (N1886, N1854, N1064, N748, N1266);
buf BUF1 (N1887, N1884);
buf BUF1 (N1888, N1871);
xor XOR2 (N1889, N1887, N523);
and AND4 (N1890, N1876, N1596, N1842, N1353);
xor XOR2 (N1891, N1873, N64);
nand NAND4 (N1892, N1889, N705, N759, N154);
buf BUF1 (N1893, N1882);
nand NAND4 (N1894, N1881, N1435, N1400, N1236);
not NOT1 (N1895, N1886);
buf BUF1 (N1896, N1892);
or OR3 (N1897, N1894, N1041, N504);
and AND4 (N1898, N1883, N370, N1830, N759);
or OR3 (N1899, N1890, N778, N899);
nor NOR3 (N1900, N1897, N1707, N263);
and AND2 (N1901, N1898, N322);
nand NAND4 (N1902, N1901, N599, N1150, N1084);
not NOT1 (N1903, N1899);
and AND4 (N1904, N1903, N630, N431, N1896);
not NOT1 (N1905, N1249);
and AND2 (N1906, N1904, N663);
nor NOR2 (N1907, N1893, N624);
and AND3 (N1908, N1879, N903, N838);
nor NOR4 (N1909, N1900, N308, N1039, N683);
xor XOR2 (N1910, N1895, N1392);
xor XOR2 (N1911, N1891, N459);
nor NOR4 (N1912, N1907, N462, N302, N1099);
nand NAND2 (N1913, N1906, N711);
not NOT1 (N1914, N1911);
xor XOR2 (N1915, N1885, N1723);
and AND4 (N1916, N1914, N435, N1081, N149);
buf BUF1 (N1917, N1908);
not NOT1 (N1918, N1888);
buf BUF1 (N1919, N1909);
nor NOR3 (N1920, N1913, N677, N59);
nand NAND3 (N1921, N1919, N1663, N95);
buf BUF1 (N1922, N1918);
and AND2 (N1923, N1922, N984);
and AND4 (N1924, N1917, N1109, N958, N453);
and AND2 (N1925, N1921, N1671);
and AND4 (N1926, N1924, N1507, N715, N1013);
or OR4 (N1927, N1910, N1632, N1403, N669);
xor XOR2 (N1928, N1916, N1264);
xor XOR2 (N1929, N1902, N1620);
and AND4 (N1930, N1929, N1569, N1453, N262);
and AND3 (N1931, N1912, N387, N1298);
and AND4 (N1932, N1915, N1784, N1465, N10);
and AND3 (N1933, N1923, N1656, N1385);
buf BUF1 (N1934, N1920);
nor NOR4 (N1935, N1930, N1007, N397, N174);
buf BUF1 (N1936, N1905);
buf BUF1 (N1937, N1928);
xor XOR2 (N1938, N1927, N1530);
not NOT1 (N1939, N1937);
and AND2 (N1940, N1932, N1769);
or OR2 (N1941, N1933, N413);
not NOT1 (N1942, N1926);
nor NOR2 (N1943, N1939, N1452);
or OR4 (N1944, N1941, N1132, N554, N351);
not NOT1 (N1945, N1943);
and AND3 (N1946, N1942, N1318, N1763);
not NOT1 (N1947, N1925);
or OR3 (N1948, N1945, N1863, N1907);
buf BUF1 (N1949, N1934);
or OR4 (N1950, N1940, N1178, N911, N1557);
nand NAND2 (N1951, N1947, N1823);
and AND4 (N1952, N1938, N79, N232, N1428);
buf BUF1 (N1953, N1935);
nor NOR4 (N1954, N1953, N635, N193, N354);
or OR4 (N1955, N1948, N191, N1304, N783);
xor XOR2 (N1956, N1952, N578);
buf BUF1 (N1957, N1944);
and AND3 (N1958, N1954, N916, N1090);
and AND3 (N1959, N1956, N1796, N1245);
and AND4 (N1960, N1949, N1925, N37, N1069);
xor XOR2 (N1961, N1951, N1334);
not NOT1 (N1962, N1931);
or OR3 (N1963, N1946, N803, N1186);
nor NOR2 (N1964, N1950, N580);
nand NAND3 (N1965, N1961, N686, N379);
and AND3 (N1966, N1964, N1587, N1529);
not NOT1 (N1967, N1963);
not NOT1 (N1968, N1957);
not NOT1 (N1969, N1967);
buf BUF1 (N1970, N1960);
nor NOR3 (N1971, N1962, N1836, N853);
xor XOR2 (N1972, N1955, N1805);
nor NOR3 (N1973, N1966, N1403, N1600);
or OR4 (N1974, N1969, N171, N1767, N1548);
xor XOR2 (N1975, N1936, N1119);
or OR4 (N1976, N1971, N994, N863, N1741);
buf BUF1 (N1977, N1973);
nor NOR2 (N1978, N1965, N1396);
or OR4 (N1979, N1968, N645, N520, N856);
buf BUF1 (N1980, N1970);
not NOT1 (N1981, N1958);
xor XOR2 (N1982, N1959, N345);
buf BUF1 (N1983, N1972);
nand NAND4 (N1984, N1979, N1933, N618, N1153);
xor XOR2 (N1985, N1978, N1053);
nand NAND3 (N1986, N1985, N1921, N143);
buf BUF1 (N1987, N1986);
not NOT1 (N1988, N1981);
xor XOR2 (N1989, N1974, N1750);
xor XOR2 (N1990, N1975, N1950);
nand NAND4 (N1991, N1977, N1778, N326, N1413);
xor XOR2 (N1992, N1987, N558);
buf BUF1 (N1993, N1988);
not NOT1 (N1994, N1983);
or OR2 (N1995, N1990, N228);
nand NAND2 (N1996, N1984, N762);
and AND4 (N1997, N1996, N390, N823, N124);
nand NAND3 (N1998, N1989, N1806, N1150);
or OR2 (N1999, N1976, N1767);
not NOT1 (N2000, N1998);
nand NAND2 (N2001, N1980, N874);
buf BUF1 (N2002, N1982);
xor XOR2 (N2003, N1995, N1964);
or OR3 (N2004, N2003, N969, N274);
xor XOR2 (N2005, N1999, N872);
nand NAND3 (N2006, N1992, N1450, N1385);
and AND4 (N2007, N2004, N1430, N1074, N338);
not NOT1 (N2008, N2006);
and AND2 (N2009, N2002, N629);
nand NAND2 (N2010, N2005, N1730);
xor XOR2 (N2011, N2008, N1294);
nor NOR2 (N2012, N2001, N1867);
and AND4 (N2013, N1994, N844, N1273, N744);
xor XOR2 (N2014, N2013, N989);
and AND4 (N2015, N2011, N572, N833, N1118);
nand NAND4 (N2016, N1993, N825, N668, N29);
and AND2 (N2017, N2012, N1553);
not NOT1 (N2018, N2007);
and AND3 (N2019, N2009, N414, N838);
nor NOR3 (N2020, N1997, N555, N499);
buf BUF1 (N2021, N2015);
xor XOR2 (N2022, N2016, N953);
not NOT1 (N2023, N2022);
and AND3 (N2024, N2014, N1079, N1684);
not NOT1 (N2025, N2023);
nor NOR3 (N2026, N2019, N1872, N913);
xor XOR2 (N2027, N2020, N1172);
nor NOR3 (N2028, N1991, N1206, N1999);
nand NAND2 (N2029, N2027, N1410);
not NOT1 (N2030, N2024);
nand NAND4 (N2031, N2018, N1826, N273, N545);
nand NAND2 (N2032, N2026, N1558);
buf BUF1 (N2033, N2030);
nand NAND4 (N2034, N2025, N862, N1666, N785);
not NOT1 (N2035, N2010);
buf BUF1 (N2036, N2029);
buf BUF1 (N2037, N2035);
nor NOR2 (N2038, N2021, N215);
not NOT1 (N2039, N2000);
nand NAND2 (N2040, N2032, N1739);
or OR3 (N2041, N2017, N372, N1936);
xor XOR2 (N2042, N2041, N689);
not NOT1 (N2043, N2039);
nand NAND3 (N2044, N2040, N717, N152);
not NOT1 (N2045, N2038);
nor NOR3 (N2046, N2037, N650, N1131);
xor XOR2 (N2047, N2046, N524);
xor XOR2 (N2048, N2043, N1946);
nor NOR4 (N2049, N2048, N300, N1143, N1484);
buf BUF1 (N2050, N2031);
buf BUF1 (N2051, N2044);
nand NAND3 (N2052, N2033, N1231, N1749);
and AND2 (N2053, N2047, N262);
xor XOR2 (N2054, N2045, N1683);
and AND2 (N2055, N2050, N267);
nand NAND2 (N2056, N2028, N349);
nor NOR4 (N2057, N2053, N208, N1286, N319);
and AND2 (N2058, N2034, N467);
or OR4 (N2059, N2055, N744, N1810, N1003);
xor XOR2 (N2060, N2049, N965);
not NOT1 (N2061, N2051);
and AND2 (N2062, N2056, N1656);
nor NOR4 (N2063, N2059, N1367, N91, N524);
and AND3 (N2064, N2060, N431, N1030);
nor NOR3 (N2065, N2042, N1474, N2026);
buf BUF1 (N2066, N2065);
or OR3 (N2067, N2057, N300, N943);
not NOT1 (N2068, N2054);
and AND4 (N2069, N2067, N1349, N231, N196);
buf BUF1 (N2070, N2036);
or OR2 (N2071, N2064, N518);
nor NOR4 (N2072, N2063, N925, N227, N1596);
buf BUF1 (N2073, N2062);
buf BUF1 (N2074, N2073);
or OR3 (N2075, N2058, N2030, N1811);
nor NOR2 (N2076, N2052, N681);
or OR3 (N2077, N2070, N977, N904);
not NOT1 (N2078, N2077);
buf BUF1 (N2079, N2072);
xor XOR2 (N2080, N2076, N1085);
nand NAND2 (N2081, N2068, N1727);
or OR3 (N2082, N2074, N1663, N487);
not NOT1 (N2083, N2082);
nand NAND4 (N2084, N2078, N1237, N211, N346);
buf BUF1 (N2085, N2066);
nor NOR4 (N2086, N2081, N573, N223, N1796);
buf BUF1 (N2087, N2071);
nand NAND3 (N2088, N2061, N1891, N1967);
nand NAND4 (N2089, N2086, N361, N1420, N471);
or OR3 (N2090, N2088, N617, N1123);
not NOT1 (N2091, N2069);
and AND2 (N2092, N2079, N18);
nand NAND2 (N2093, N2090, N575);
nand NAND4 (N2094, N2084, N238, N1520, N1720);
and AND4 (N2095, N2091, N1068, N849, N1574);
xor XOR2 (N2096, N2095, N1592);
buf BUF1 (N2097, N2083);
nor NOR2 (N2098, N2094, N614);
not NOT1 (N2099, N2096);
not NOT1 (N2100, N2097);
not NOT1 (N2101, N2075);
xor XOR2 (N2102, N2101, N1840);
buf BUF1 (N2103, N2087);
nand NAND3 (N2104, N2080, N141, N1654);
buf BUF1 (N2105, N2102);
nand NAND3 (N2106, N2085, N2104, N1066);
xor XOR2 (N2107, N509, N1999);
not NOT1 (N2108, N2105);
nand NAND2 (N2109, N2100, N1235);
nand NAND4 (N2110, N2089, N1785, N2012, N252);
xor XOR2 (N2111, N2110, N2009);
and AND3 (N2112, N2098, N1770, N1952);
and AND2 (N2113, N2093, N695);
and AND2 (N2114, N2092, N96);
nor NOR4 (N2115, N2114, N768, N406, N1012);
or OR3 (N2116, N2109, N294, N794);
nor NOR3 (N2117, N2115, N1077, N1166);
buf BUF1 (N2118, N2111);
nor NOR2 (N2119, N2106, N1492);
or OR4 (N2120, N2118, N1855, N1545, N1369);
nand NAND4 (N2121, N2103, N44, N1281, N1248);
xor XOR2 (N2122, N2119, N1815);
nor NOR2 (N2123, N2108, N1667);
buf BUF1 (N2124, N2113);
not NOT1 (N2125, N2116);
xor XOR2 (N2126, N2122, N850);
or OR3 (N2127, N2124, N1159, N1651);
not NOT1 (N2128, N2126);
or OR3 (N2129, N2127, N1630, N509);
nand NAND3 (N2130, N2123, N577, N465);
and AND3 (N2131, N2120, N774, N1166);
not NOT1 (N2132, N2130);
and AND3 (N2133, N2117, N264, N1745);
xor XOR2 (N2134, N2133, N610);
and AND3 (N2135, N2125, N1832, N247);
buf BUF1 (N2136, N2128);
buf BUF1 (N2137, N2129);
or OR3 (N2138, N2131, N760, N545);
and AND4 (N2139, N2138, N410, N791, N1383);
or OR2 (N2140, N2132, N796);
not NOT1 (N2141, N2140);
xor XOR2 (N2142, N2141, N1325);
nor NOR2 (N2143, N2121, N1342);
nor NOR3 (N2144, N2142, N28, N749);
buf BUF1 (N2145, N2139);
not NOT1 (N2146, N2099);
nand NAND2 (N2147, N2134, N2056);
and AND4 (N2148, N2137, N1398, N566, N1503);
buf BUF1 (N2149, N2147);
nand NAND3 (N2150, N2112, N755, N1024);
or OR2 (N2151, N2144, N1167);
buf BUF1 (N2152, N2107);
buf BUF1 (N2153, N2146);
buf BUF1 (N2154, N2153);
nor NOR3 (N2155, N2151, N1934, N1472);
or OR3 (N2156, N2149, N1898, N1658);
xor XOR2 (N2157, N2156, N183);
nand NAND2 (N2158, N2136, N593);
or OR4 (N2159, N2150, N1846, N2147, N2138);
nor NOR2 (N2160, N2154, N1329);
or OR3 (N2161, N2148, N1900, N805);
or OR2 (N2162, N2159, N1315);
buf BUF1 (N2163, N2161);
nand NAND4 (N2164, N2135, N34, N126, N958);
or OR4 (N2165, N2157, N1348, N407, N1021);
nor NOR3 (N2166, N2152, N2116, N1054);
buf BUF1 (N2167, N2166);
not NOT1 (N2168, N2163);
buf BUF1 (N2169, N2167);
not NOT1 (N2170, N2158);
buf BUF1 (N2171, N2169);
nand NAND4 (N2172, N2165, N1560, N1197, N1145);
xor XOR2 (N2173, N2171, N1002);
nor NOR2 (N2174, N2160, N1363);
nand NAND4 (N2175, N2170, N478, N1655, N621);
xor XOR2 (N2176, N2175, N2099);
nor NOR3 (N2177, N2168, N42, N2052);
not NOT1 (N2178, N2164);
not NOT1 (N2179, N2178);
xor XOR2 (N2180, N2155, N296);
nor NOR2 (N2181, N2179, N2079);
not NOT1 (N2182, N2174);
or OR2 (N2183, N2182, N156);
buf BUF1 (N2184, N2180);
xor XOR2 (N2185, N2177, N1676);
nand NAND2 (N2186, N2181, N17);
nor NOR3 (N2187, N2176, N1089, N1886);
or OR2 (N2188, N2185, N621);
nand NAND4 (N2189, N2187, N1279, N618, N1924);
xor XOR2 (N2190, N2162, N1350);
and AND4 (N2191, N2188, N1609, N1396, N258);
xor XOR2 (N2192, N2184, N347);
or OR4 (N2193, N2173, N582, N981, N1489);
nand NAND2 (N2194, N2145, N1499);
buf BUF1 (N2195, N2194);
not NOT1 (N2196, N2183);
not NOT1 (N2197, N2196);
nor NOR2 (N2198, N2190, N2071);
not NOT1 (N2199, N2195);
not NOT1 (N2200, N2198);
nand NAND2 (N2201, N2192, N1375);
and AND3 (N2202, N2143, N322, N1138);
or OR3 (N2203, N2193, N1979, N2175);
not NOT1 (N2204, N2201);
not NOT1 (N2205, N2202);
nand NAND3 (N2206, N2197, N354, N1670);
not NOT1 (N2207, N2206);
nor NOR2 (N2208, N2205, N2140);
not NOT1 (N2209, N2208);
nor NOR4 (N2210, N2199, N1419, N1650, N1404);
nand NAND4 (N2211, N2204, N1602, N184, N1322);
nor NOR2 (N2212, N2211, N991);
xor XOR2 (N2213, N2203, N1949);
nand NAND4 (N2214, N2207, N1403, N51, N2194);
or OR4 (N2215, N2209, N163, N130, N2148);
nor NOR2 (N2216, N2189, N2132);
and AND2 (N2217, N2216, N1333);
or OR3 (N2218, N2186, N946, N1916);
not NOT1 (N2219, N2200);
buf BUF1 (N2220, N2191);
nand NAND2 (N2221, N2217, N686);
and AND2 (N2222, N2221, N603);
nor NOR2 (N2223, N2210, N409);
not NOT1 (N2224, N2220);
not NOT1 (N2225, N2219);
buf BUF1 (N2226, N2213);
nor NOR4 (N2227, N2172, N136, N44, N1113);
nor NOR3 (N2228, N2222, N908, N67);
and AND2 (N2229, N2212, N877);
xor XOR2 (N2230, N2225, N78);
not NOT1 (N2231, N2227);
buf BUF1 (N2232, N2231);
nor NOR4 (N2233, N2226, N952, N1983, N863);
nor NOR4 (N2234, N2232, N985, N1588, N1231);
buf BUF1 (N2235, N2215);
and AND2 (N2236, N2214, N1246);
buf BUF1 (N2237, N2229);
xor XOR2 (N2238, N2236, N704);
nand NAND2 (N2239, N2218, N1846);
xor XOR2 (N2240, N2233, N734);
buf BUF1 (N2241, N2239);
buf BUF1 (N2242, N2241);
nor NOR3 (N2243, N2230, N115, N501);
nand NAND2 (N2244, N2242, N111);
nor NOR4 (N2245, N2224, N1769, N1652, N353);
xor XOR2 (N2246, N2238, N629);
and AND3 (N2247, N2246, N999, N1185);
nor NOR4 (N2248, N2243, N344, N1776, N1020);
not NOT1 (N2249, N2223);
nand NAND2 (N2250, N2235, N1257);
buf BUF1 (N2251, N2237);
nor NOR3 (N2252, N2248, N404, N464);
and AND3 (N2253, N2240, N716, N113);
and AND3 (N2254, N2250, N468, N873);
nand NAND2 (N2255, N2251, N122);
nand NAND2 (N2256, N2228, N257);
or OR4 (N2257, N2234, N899, N1256, N2187);
nor NOR2 (N2258, N2256, N1698);
and AND4 (N2259, N2255, N1275, N1298, N2236);
or OR3 (N2260, N2244, N718, N133);
buf BUF1 (N2261, N2257);
buf BUF1 (N2262, N2260);
nor NOR3 (N2263, N2245, N1761, N1949);
not NOT1 (N2264, N2263);
and AND3 (N2265, N2252, N1925, N317);
nor NOR4 (N2266, N2261, N228, N360, N1352);
nor NOR2 (N2267, N2254, N1227);
nand NAND3 (N2268, N2253, N1470, N1192);
and AND3 (N2269, N2258, N921, N505);
or OR4 (N2270, N2268, N574, N119, N1137);
not NOT1 (N2271, N2264);
buf BUF1 (N2272, N2247);
nand NAND3 (N2273, N2271, N1208, N1367);
and AND3 (N2274, N2267, N2179, N2023);
buf BUF1 (N2275, N2272);
buf BUF1 (N2276, N2273);
xor XOR2 (N2277, N2266, N1394);
buf BUF1 (N2278, N2265);
nor NOR4 (N2279, N2276, N1548, N1203, N1166);
and AND2 (N2280, N2275, N1363);
xor XOR2 (N2281, N2249, N1702);
nand NAND4 (N2282, N2270, N1816, N418, N1830);
or OR4 (N2283, N2277, N2002, N757, N793);
buf BUF1 (N2284, N2278);
not NOT1 (N2285, N2274);
nor NOR2 (N2286, N2280, N1847);
and AND3 (N2287, N2281, N656, N1226);
buf BUF1 (N2288, N2259);
not NOT1 (N2289, N2287);
not NOT1 (N2290, N2282);
not NOT1 (N2291, N2283);
or OR2 (N2292, N2289, N402);
nand NAND3 (N2293, N2269, N1064, N2201);
xor XOR2 (N2294, N2285, N749);
nand NAND2 (N2295, N2279, N1249);
and AND2 (N2296, N2295, N130);
not NOT1 (N2297, N2286);
nand NAND3 (N2298, N2290, N144, N1265);
not NOT1 (N2299, N2294);
buf BUF1 (N2300, N2284);
nor NOR4 (N2301, N2296, N1091, N181, N888);
and AND2 (N2302, N2298, N113);
xor XOR2 (N2303, N2297, N810);
buf BUF1 (N2304, N2300);
buf BUF1 (N2305, N2303);
nand NAND3 (N2306, N2292, N2070, N613);
and AND4 (N2307, N2291, N151, N1947, N1600);
and AND2 (N2308, N2302, N1662);
or OR4 (N2309, N2288, N243, N1713, N2060);
and AND4 (N2310, N2262, N1554, N1362, N131);
buf BUF1 (N2311, N2304);
nor NOR4 (N2312, N2299, N847, N1936, N2106);
buf BUF1 (N2313, N2293);
nor NOR2 (N2314, N2310, N2031);
not NOT1 (N2315, N2301);
nor NOR2 (N2316, N2314, N1230);
not NOT1 (N2317, N2311);
and AND4 (N2318, N2316, N699, N873, N468);
buf BUF1 (N2319, N2305);
nand NAND2 (N2320, N2309, N1876);
buf BUF1 (N2321, N2312);
nand NAND3 (N2322, N2307, N1256, N1576);
or OR3 (N2323, N2306, N1978, N174);
and AND4 (N2324, N2313, N2052, N1884, N45);
or OR2 (N2325, N2324, N1653);
nand NAND4 (N2326, N2317, N293, N1087, N1671);
not NOT1 (N2327, N2322);
and AND4 (N2328, N2320, N1483, N1534, N1900);
or OR2 (N2329, N2326, N1817);
and AND3 (N2330, N2329, N445, N61);
nor NOR4 (N2331, N2325, N1912, N1478, N2040);
buf BUF1 (N2332, N2328);
or OR4 (N2333, N2323, N1745, N1947, N2125);
xor XOR2 (N2334, N2315, N872);
nor NOR2 (N2335, N2334, N1459);
buf BUF1 (N2336, N2308);
and AND4 (N2337, N2319, N1794, N2212, N559);
nor NOR2 (N2338, N2335, N1354);
buf BUF1 (N2339, N2337);
and AND2 (N2340, N2336, N123);
xor XOR2 (N2341, N2318, N1263);
not NOT1 (N2342, N2339);
buf BUF1 (N2343, N2340);
buf BUF1 (N2344, N2338);
nand NAND4 (N2345, N2343, N1373, N807, N2022);
buf BUF1 (N2346, N2321);
xor XOR2 (N2347, N2344, N886);
or OR2 (N2348, N2346, N621);
nand NAND3 (N2349, N2333, N615, N1815);
not NOT1 (N2350, N2349);
buf BUF1 (N2351, N2327);
nor NOR4 (N2352, N2341, N186, N1835, N51);
buf BUF1 (N2353, N2347);
nand NAND4 (N2354, N2331, N876, N1446, N875);
xor XOR2 (N2355, N2353, N2013);
nor NOR2 (N2356, N2345, N2005);
xor XOR2 (N2357, N2351, N332);
buf BUF1 (N2358, N2332);
nor NOR4 (N2359, N2342, N1215, N2144, N1019);
buf BUF1 (N2360, N2350);
buf BUF1 (N2361, N2357);
buf BUF1 (N2362, N2348);
or OR4 (N2363, N2352, N874, N1312, N824);
nand NAND3 (N2364, N2363, N1431, N477);
not NOT1 (N2365, N2356);
nor NOR4 (N2366, N2354, N1337, N1842, N548);
not NOT1 (N2367, N2359);
nor NOR3 (N2368, N2355, N133, N2055);
not NOT1 (N2369, N2360);
xor XOR2 (N2370, N2368, N1859);
and AND2 (N2371, N2362, N2266);
or OR2 (N2372, N2371, N1743);
xor XOR2 (N2373, N2366, N2369);
not NOT1 (N2374, N1325);
not NOT1 (N2375, N2364);
nand NAND2 (N2376, N2358, N1765);
not NOT1 (N2377, N2373);
or OR2 (N2378, N2375, N610);
xor XOR2 (N2379, N2370, N1874);
not NOT1 (N2380, N2374);
not NOT1 (N2381, N2379);
buf BUF1 (N2382, N2367);
and AND4 (N2383, N2380, N493, N1342, N1560);
not NOT1 (N2384, N2382);
xor XOR2 (N2385, N2378, N2010);
nand NAND3 (N2386, N2377, N2087, N1638);
xor XOR2 (N2387, N2365, N23);
not NOT1 (N2388, N2361);
and AND3 (N2389, N2376, N1344, N78);
nand NAND2 (N2390, N2388, N982);
nand NAND4 (N2391, N2385, N937, N1724, N104);
or OR4 (N2392, N2381, N1282, N2066, N338);
nand NAND3 (N2393, N2330, N1710, N1439);
nand NAND2 (N2394, N2391, N1826);
or OR3 (N2395, N2383, N2307, N1394);
not NOT1 (N2396, N2387);
and AND4 (N2397, N2392, N1122, N198, N456);
nand NAND2 (N2398, N2390, N933);
nand NAND2 (N2399, N2384, N596);
not NOT1 (N2400, N2397);
not NOT1 (N2401, N2386);
xor XOR2 (N2402, N2400, N676);
xor XOR2 (N2403, N2394, N1733);
nor NOR3 (N2404, N2372, N1652, N2342);
not NOT1 (N2405, N2399);
nor NOR4 (N2406, N2402, N147, N1045, N2223);
not NOT1 (N2407, N2405);
buf BUF1 (N2408, N2404);
buf BUF1 (N2409, N2395);
and AND2 (N2410, N2403, N1169);
and AND4 (N2411, N2393, N2185, N2041, N1307);
buf BUF1 (N2412, N2411);
or OR4 (N2413, N2401, N1168, N1205, N476);
nor NOR2 (N2414, N2412, N2166);
nor NOR2 (N2415, N2407, N1370);
or OR4 (N2416, N2406, N336, N1833, N1894);
xor XOR2 (N2417, N2409, N2005);
or OR2 (N2418, N2415, N1149);
xor XOR2 (N2419, N2396, N641);
and AND2 (N2420, N2408, N2163);
nand NAND4 (N2421, N2398, N1429, N305, N798);
and AND4 (N2422, N2418, N1196, N1028, N495);
nand NAND2 (N2423, N2416, N963);
not NOT1 (N2424, N2420);
or OR3 (N2425, N2389, N934, N1454);
or OR3 (N2426, N2413, N2007, N2129);
nor NOR2 (N2427, N2425, N2041);
not NOT1 (N2428, N2410);
nor NOR2 (N2429, N2414, N1575);
nand NAND2 (N2430, N2423, N460);
or OR2 (N2431, N2424, N357);
buf BUF1 (N2432, N2427);
xor XOR2 (N2433, N2419, N697);
and AND3 (N2434, N2428, N1227, N1709);
xor XOR2 (N2435, N2421, N1902);
not NOT1 (N2436, N2422);
not NOT1 (N2437, N2433);
xor XOR2 (N2438, N2431, N848);
xor XOR2 (N2439, N2437, N1283);
nor NOR3 (N2440, N2430, N394, N1272);
nor NOR4 (N2441, N2435, N979, N2310, N1756);
xor XOR2 (N2442, N2436, N2069);
nor NOR3 (N2443, N2426, N84, N1270);
buf BUF1 (N2444, N2443);
xor XOR2 (N2445, N2434, N76);
nor NOR3 (N2446, N2445, N1541, N887);
and AND3 (N2447, N2429, N1550, N1786);
nor NOR3 (N2448, N2440, N2048, N2105);
xor XOR2 (N2449, N2442, N1042);
not NOT1 (N2450, N2438);
and AND3 (N2451, N2444, N1101, N1524);
and AND3 (N2452, N2432, N198, N478);
xor XOR2 (N2453, N2439, N871);
xor XOR2 (N2454, N2448, N1036);
nand NAND2 (N2455, N2453, N75);
xor XOR2 (N2456, N2451, N1951);
nor NOR4 (N2457, N2452, N1995, N1329, N1288);
xor XOR2 (N2458, N2447, N2288);
buf BUF1 (N2459, N2457);
nand NAND4 (N2460, N2449, N1367, N1632, N1412);
not NOT1 (N2461, N2441);
xor XOR2 (N2462, N2460, N1761);
or OR3 (N2463, N2458, N2003, N688);
buf BUF1 (N2464, N2446);
nand NAND2 (N2465, N2464, N305);
xor XOR2 (N2466, N2417, N1039);
not NOT1 (N2467, N2454);
xor XOR2 (N2468, N2450, N544);
nand NAND2 (N2469, N2459, N1002);
nor NOR2 (N2470, N2461, N892);
and AND3 (N2471, N2468, N1652, N2176);
not NOT1 (N2472, N2471);
xor XOR2 (N2473, N2465, N1243);
nor NOR3 (N2474, N2466, N1954, N1538);
buf BUF1 (N2475, N2473);
or OR4 (N2476, N2474, N737, N1207, N1936);
not NOT1 (N2477, N2475);
xor XOR2 (N2478, N2462, N2246);
and AND4 (N2479, N2455, N2072, N613, N149);
nor NOR3 (N2480, N2477, N609, N1586);
or OR3 (N2481, N2470, N329, N2290);
not NOT1 (N2482, N2479);
or OR3 (N2483, N2472, N200, N1690);
and AND4 (N2484, N2481, N305, N1503, N1133);
xor XOR2 (N2485, N2484, N105);
buf BUF1 (N2486, N2483);
buf BUF1 (N2487, N2467);
not NOT1 (N2488, N2469);
nor NOR3 (N2489, N2485, N268, N2298);
nor NOR2 (N2490, N2456, N2316);
nand NAND3 (N2491, N2463, N63, N1458);
not NOT1 (N2492, N2487);
xor XOR2 (N2493, N2488, N1152);
buf BUF1 (N2494, N2486);
xor XOR2 (N2495, N2493, N1437);
buf BUF1 (N2496, N2489);
nand NAND4 (N2497, N2490, N13, N1991, N684);
buf BUF1 (N2498, N2494);
nand NAND4 (N2499, N2495, N538, N295, N896);
buf BUF1 (N2500, N2497);
xor XOR2 (N2501, N2491, N1022);
and AND2 (N2502, N2501, N2057);
or OR3 (N2503, N2482, N159, N1478);
nand NAND3 (N2504, N2500, N1612, N604);
buf BUF1 (N2505, N2478);
nand NAND4 (N2506, N2492, N53, N332, N2403);
nor NOR3 (N2507, N2476, N900, N463);
or OR2 (N2508, N2504, N1970);
xor XOR2 (N2509, N2496, N657);
and AND4 (N2510, N2480, N232, N594, N2183);
nand NAND4 (N2511, N2503, N2418, N1219, N315);
xor XOR2 (N2512, N2498, N138);
and AND4 (N2513, N2510, N1845, N980, N896);
xor XOR2 (N2514, N2511, N2365);
nand NAND2 (N2515, N2514, N1299);
buf BUF1 (N2516, N2515);
and AND4 (N2517, N2507, N1554, N771, N266);
not NOT1 (N2518, N2502);
buf BUF1 (N2519, N2518);
nand NAND4 (N2520, N2517, N1040, N1163, N2092);
xor XOR2 (N2521, N2499, N925);
not NOT1 (N2522, N2508);
buf BUF1 (N2523, N2505);
buf BUF1 (N2524, N2521);
not NOT1 (N2525, N2520);
nor NOR2 (N2526, N2519, N1822);
or OR2 (N2527, N2506, N50);
and AND4 (N2528, N2522, N930, N857, N1556);
and AND4 (N2529, N2524, N1661, N1694, N2306);
xor XOR2 (N2530, N2513, N742);
nand NAND3 (N2531, N2525, N2415, N873);
and AND4 (N2532, N2512, N1072, N507, N2168);
buf BUF1 (N2533, N2532);
or OR4 (N2534, N2509, N435, N988, N1764);
nor NOR4 (N2535, N2516, N1136, N1649, N639);
not NOT1 (N2536, N2531);
nor NOR4 (N2537, N2528, N479, N1210, N2447);
nor NOR3 (N2538, N2534, N750, N2106);
or OR2 (N2539, N2535, N239);
nand NAND2 (N2540, N2529, N1565);
buf BUF1 (N2541, N2523);
xor XOR2 (N2542, N2538, N661);
nor NOR2 (N2543, N2527, N300);
not NOT1 (N2544, N2542);
nand NAND2 (N2545, N2541, N1736);
or OR3 (N2546, N2536, N1074, N1715);
or OR4 (N2547, N2539, N1308, N1600, N665);
nand NAND2 (N2548, N2540, N2533);
nor NOR4 (N2549, N604, N2358, N2270, N1310);
and AND3 (N2550, N2537, N87, N430);
or OR4 (N2551, N2543, N2489, N218, N585);
or OR3 (N2552, N2545, N876, N977);
buf BUF1 (N2553, N2551);
buf BUF1 (N2554, N2550);
xor XOR2 (N2555, N2530, N1898);
not NOT1 (N2556, N2526);
and AND2 (N2557, N2554, N1542);
not NOT1 (N2558, N2544);
nand NAND4 (N2559, N2549, N542, N1922, N1052);
xor XOR2 (N2560, N2559, N833);
and AND3 (N2561, N2557, N1183, N852);
or OR3 (N2562, N2552, N61, N2200);
buf BUF1 (N2563, N2553);
xor XOR2 (N2564, N2560, N2104);
not NOT1 (N2565, N2555);
not NOT1 (N2566, N2565);
buf BUF1 (N2567, N2546);
xor XOR2 (N2568, N2556, N1946);
xor XOR2 (N2569, N2566, N1875);
nand NAND3 (N2570, N2568, N1282, N2026);
or OR4 (N2571, N2548, N2301, N2428, N664);
not NOT1 (N2572, N2571);
or OR4 (N2573, N2564, N449, N2300, N63);
buf BUF1 (N2574, N2567);
xor XOR2 (N2575, N2547, N941);
xor XOR2 (N2576, N2562, N2301);
nor NOR2 (N2577, N2558, N2344);
not NOT1 (N2578, N2574);
buf BUF1 (N2579, N2561);
and AND3 (N2580, N2579, N1478, N601);
xor XOR2 (N2581, N2576, N1471);
xor XOR2 (N2582, N2573, N921);
and AND3 (N2583, N2582, N255, N789);
not NOT1 (N2584, N2563);
xor XOR2 (N2585, N2572, N208);
and AND4 (N2586, N2575, N473, N1240, N1910);
xor XOR2 (N2587, N2583, N1891);
buf BUF1 (N2588, N2585);
nand NAND3 (N2589, N2569, N146, N705);
not NOT1 (N2590, N2577);
not NOT1 (N2591, N2581);
and AND3 (N2592, N2578, N2306, N28);
or OR3 (N2593, N2587, N1804, N2161);
buf BUF1 (N2594, N2593);
xor XOR2 (N2595, N2591, N2028);
and AND4 (N2596, N2594, N2052, N1536, N2258);
not NOT1 (N2597, N2596);
or OR3 (N2598, N2590, N11, N501);
nor NOR2 (N2599, N2586, N962);
and AND2 (N2600, N2595, N1870);
nor NOR2 (N2601, N2589, N2084);
or OR3 (N2602, N2597, N2258, N1688);
xor XOR2 (N2603, N2600, N2128);
buf BUF1 (N2604, N2602);
not NOT1 (N2605, N2604);
xor XOR2 (N2606, N2592, N2291);
or OR2 (N2607, N2605, N1878);
and AND4 (N2608, N2588, N845, N1824, N2108);
not NOT1 (N2609, N2608);
nand NAND4 (N2610, N2609, N206, N1073, N1583);
nand NAND4 (N2611, N2606, N277, N2411, N2132);
not NOT1 (N2612, N2584);
or OR4 (N2613, N2610, N2041, N1529, N1684);
not NOT1 (N2614, N2598);
xor XOR2 (N2615, N2570, N2089);
and AND2 (N2616, N2614, N1476);
nor NOR4 (N2617, N2611, N1510, N790, N1251);
buf BUF1 (N2618, N2616);
and AND3 (N2619, N2601, N507, N666);
and AND3 (N2620, N2580, N1226, N2544);
not NOT1 (N2621, N2613);
nor NOR4 (N2622, N2618, N2023, N1101, N491);
and AND3 (N2623, N2612, N1448, N2343);
xor XOR2 (N2624, N2607, N465);
and AND3 (N2625, N2624, N796, N2079);
nand NAND4 (N2626, N2599, N1755, N2295, N2137);
xor XOR2 (N2627, N2621, N1194);
nand NAND3 (N2628, N2619, N2463, N779);
not NOT1 (N2629, N2626);
or OR2 (N2630, N2603, N1426);
or OR2 (N2631, N2629, N2616);
nor NOR4 (N2632, N2617, N1540, N1466, N389);
or OR4 (N2633, N2630, N1278, N1423, N309);
and AND4 (N2634, N2625, N891, N1012, N2005);
xor XOR2 (N2635, N2633, N82);
or OR3 (N2636, N2620, N637, N1195);
nand NAND4 (N2637, N2627, N257, N712, N1128);
buf BUF1 (N2638, N2631);
xor XOR2 (N2639, N2636, N1990);
xor XOR2 (N2640, N2632, N1294);
buf BUF1 (N2641, N2635);
xor XOR2 (N2642, N2615, N1381);
not NOT1 (N2643, N2638);
not NOT1 (N2644, N2642);
buf BUF1 (N2645, N2623);
buf BUF1 (N2646, N2640);
and AND4 (N2647, N2628, N2074, N1115, N1776);
not NOT1 (N2648, N2634);
nor NOR2 (N2649, N2647, N147);
and AND2 (N2650, N2646, N675);
xor XOR2 (N2651, N2650, N2329);
nor NOR4 (N2652, N2649, N958, N1064, N2163);
and AND4 (N2653, N2645, N2487, N2019, N1661);
nand NAND4 (N2654, N2652, N1623, N1957, N1612);
buf BUF1 (N2655, N2648);
not NOT1 (N2656, N2622);
or OR2 (N2657, N2641, N983);
not NOT1 (N2658, N2654);
nand NAND3 (N2659, N2639, N177, N2348);
xor XOR2 (N2660, N2655, N1807);
and AND4 (N2661, N2637, N1961, N694, N48);
nor NOR4 (N2662, N2644, N1721, N1483, N1305);
buf BUF1 (N2663, N2661);
or OR3 (N2664, N2660, N312, N922);
buf BUF1 (N2665, N2664);
or OR2 (N2666, N2651, N1027);
nand NAND2 (N2667, N2665, N775);
not NOT1 (N2668, N2662);
buf BUF1 (N2669, N2658);
not NOT1 (N2670, N2668);
or OR3 (N2671, N2659, N1944, N521);
or OR4 (N2672, N2671, N2382, N1244, N841);
or OR3 (N2673, N2669, N1704, N994);
buf BUF1 (N2674, N2653);
and AND3 (N2675, N2674, N1983, N2091);
and AND3 (N2676, N2643, N885, N1323);
buf BUF1 (N2677, N2666);
buf BUF1 (N2678, N2676);
nand NAND3 (N2679, N2656, N2485, N1606);
xor XOR2 (N2680, N2678, N2644);
or OR4 (N2681, N2657, N2512, N2084, N2397);
xor XOR2 (N2682, N2667, N2368);
or OR2 (N2683, N2682, N623);
buf BUF1 (N2684, N2675);
nand NAND4 (N2685, N2680, N1993, N2486, N1932);
nor NOR2 (N2686, N2677, N1650);
and AND2 (N2687, N2684, N714);
buf BUF1 (N2688, N2683);
or OR4 (N2689, N2670, N757, N699, N417);
buf BUF1 (N2690, N2686);
or OR2 (N2691, N2672, N86);
nand NAND3 (N2692, N2690, N414, N581);
nor NOR3 (N2693, N2689, N2044, N2145);
nand NAND4 (N2694, N2673, N1522, N2369, N132);
xor XOR2 (N2695, N2688, N1176);
nor NOR3 (N2696, N2692, N1915, N769);
buf BUF1 (N2697, N2681);
nand NAND4 (N2698, N2693, N1942, N22, N1367);
buf BUF1 (N2699, N2663);
not NOT1 (N2700, N2696);
and AND2 (N2701, N2699, N1707);
nor NOR3 (N2702, N2679, N51, N524);
nand NAND3 (N2703, N2685, N2366, N962);
and AND3 (N2704, N2702, N619, N2011);
nor NOR2 (N2705, N2700, N709);
not NOT1 (N2706, N2697);
nand NAND2 (N2707, N2703, N965);
xor XOR2 (N2708, N2701, N932);
nand NAND4 (N2709, N2705, N2659, N1002, N924);
nand NAND2 (N2710, N2707, N850);
xor XOR2 (N2711, N2694, N2544);
not NOT1 (N2712, N2710);
nand NAND2 (N2713, N2708, N2203);
and AND3 (N2714, N2698, N1754, N1000);
not NOT1 (N2715, N2687);
or OR3 (N2716, N2709, N1019, N2195);
xor XOR2 (N2717, N2711, N445);
or OR4 (N2718, N2716, N2299, N657, N1659);
nor NOR3 (N2719, N2695, N959, N1752);
xor XOR2 (N2720, N2719, N373);
buf BUF1 (N2721, N2691);
xor XOR2 (N2722, N2720, N2307);
nor NOR3 (N2723, N2712, N2177, N400);
buf BUF1 (N2724, N2723);
and AND4 (N2725, N2714, N2358, N2330, N1164);
xor XOR2 (N2726, N2715, N249);
and AND4 (N2727, N2713, N831, N684, N1899);
or OR4 (N2728, N2722, N2584, N1460, N2439);
not NOT1 (N2729, N2727);
xor XOR2 (N2730, N2726, N2133);
or OR2 (N2731, N2721, N2035);
xor XOR2 (N2732, N2730, N448);
and AND3 (N2733, N2724, N2405, N1298);
or OR3 (N2734, N2725, N332, N2001);
nor NOR2 (N2735, N2734, N1222);
and AND4 (N2736, N2733, N1116, N67, N423);
nor NOR2 (N2737, N2732, N2228);
xor XOR2 (N2738, N2717, N161);
xor XOR2 (N2739, N2738, N35);
xor XOR2 (N2740, N2736, N1565);
nor NOR2 (N2741, N2740, N798);
nand NAND3 (N2742, N2718, N2135, N1052);
and AND3 (N2743, N2731, N1627, N2450);
nand NAND4 (N2744, N2743, N360, N417, N2067);
or OR4 (N2745, N2704, N2369, N866, N1962);
not NOT1 (N2746, N2729);
not NOT1 (N2747, N2741);
buf BUF1 (N2748, N2737);
not NOT1 (N2749, N2739);
nand NAND4 (N2750, N2735, N1914, N2478, N2343);
buf BUF1 (N2751, N2728);
nor NOR2 (N2752, N2745, N572);
nor NOR3 (N2753, N2751, N1188, N1988);
nor NOR4 (N2754, N2742, N1252, N255, N1549);
not NOT1 (N2755, N2748);
or OR3 (N2756, N2750, N2024, N570);
xor XOR2 (N2757, N2749, N1345);
xor XOR2 (N2758, N2754, N696);
or OR2 (N2759, N2747, N2252);
not NOT1 (N2760, N2759);
nor NOR2 (N2761, N2756, N630);
xor XOR2 (N2762, N2746, N210);
nor NOR2 (N2763, N2744, N1422);
xor XOR2 (N2764, N2757, N397);
and AND3 (N2765, N2752, N765, N732);
or OR2 (N2766, N2706, N1503);
nand NAND4 (N2767, N2764, N584, N2268, N1829);
xor XOR2 (N2768, N2762, N1277);
or OR2 (N2769, N2765, N2766);
xor XOR2 (N2770, N262, N2011);
not NOT1 (N2771, N2755);
not NOT1 (N2772, N2771);
buf BUF1 (N2773, N2763);
or OR2 (N2774, N2772, N725);
buf BUF1 (N2775, N2769);
not NOT1 (N2776, N2758);
not NOT1 (N2777, N2770);
or OR4 (N2778, N2761, N1163, N2163, N1708);
not NOT1 (N2779, N2776);
buf BUF1 (N2780, N2768);
nand NAND3 (N2781, N2760, N2738, N2255);
nand NAND2 (N2782, N2779, N2230);
or OR2 (N2783, N2774, N2223);
nor NOR3 (N2784, N2753, N1096, N1340);
not NOT1 (N2785, N2783);
nor NOR2 (N2786, N2781, N2045);
nand NAND2 (N2787, N2782, N2249);
and AND4 (N2788, N2786, N782, N2515, N2492);
or OR4 (N2789, N2785, N788, N1480, N104);
not NOT1 (N2790, N2773);
and AND2 (N2791, N2790, N409);
nand NAND4 (N2792, N2784, N1244, N1577, N1991);
or OR4 (N2793, N2789, N225, N1517, N1602);
not NOT1 (N2794, N2788);
and AND2 (N2795, N2792, N1125);
buf BUF1 (N2796, N2777);
not NOT1 (N2797, N2794);
and AND4 (N2798, N2787, N1026, N1583, N1482);
not NOT1 (N2799, N2798);
or OR4 (N2800, N2795, N2519, N1535, N118);
buf BUF1 (N2801, N2799);
nand NAND4 (N2802, N2778, N2743, N350, N671);
buf BUF1 (N2803, N2791);
buf BUF1 (N2804, N2780);
nor NOR2 (N2805, N2802, N2750);
nor NOR2 (N2806, N2775, N2226);
or OR2 (N2807, N2805, N786);
nor NOR3 (N2808, N2806, N1401, N2422);
and AND3 (N2809, N2767, N1612, N1720);
nor NOR2 (N2810, N2800, N1374);
not NOT1 (N2811, N2797);
xor XOR2 (N2812, N2803, N2454);
nand NAND2 (N2813, N2810, N412);
xor XOR2 (N2814, N2812, N2154);
and AND3 (N2815, N2801, N113, N139);
and AND3 (N2816, N2813, N1274, N912);
buf BUF1 (N2817, N2804);
and AND2 (N2818, N2808, N162);
nand NAND3 (N2819, N2816, N684, N941);
or OR2 (N2820, N2811, N1717);
xor XOR2 (N2821, N2817, N1926);
buf BUF1 (N2822, N2809);
or OR2 (N2823, N2807, N2690);
or OR4 (N2824, N2823, N1446, N1107, N2641);
nor NOR3 (N2825, N2819, N49, N1646);
xor XOR2 (N2826, N2793, N1030);
or OR3 (N2827, N2826, N210, N1198);
nor NOR2 (N2828, N2814, N2755);
buf BUF1 (N2829, N2822);
xor XOR2 (N2830, N2818, N2085);
and AND4 (N2831, N2796, N2107, N2699, N1755);
buf BUF1 (N2832, N2820);
not NOT1 (N2833, N2815);
buf BUF1 (N2834, N2830);
xor XOR2 (N2835, N2827, N1702);
nor NOR3 (N2836, N2831, N2188, N2329);
or OR3 (N2837, N2835, N133, N980);
and AND4 (N2838, N2828, N1460, N346, N2269);
and AND4 (N2839, N2821, N1896, N685, N1790);
buf BUF1 (N2840, N2833);
and AND3 (N2841, N2839, N1920, N2216);
buf BUF1 (N2842, N2825);
nand NAND3 (N2843, N2834, N132, N1253);
or OR3 (N2844, N2832, N2654, N1151);
and AND3 (N2845, N2837, N1323, N1709);
and AND4 (N2846, N2843, N1163, N2303, N1835);
not NOT1 (N2847, N2842);
or OR2 (N2848, N2847, N518);
nand NAND4 (N2849, N2824, N1355, N100, N973);
or OR2 (N2850, N2838, N603);
xor XOR2 (N2851, N2844, N61);
nor NOR2 (N2852, N2840, N2108);
nor NOR2 (N2853, N2841, N2379);
nand NAND3 (N2854, N2836, N1244, N2571);
nand NAND3 (N2855, N2851, N1316, N1116);
xor XOR2 (N2856, N2829, N2546);
not NOT1 (N2857, N2853);
or OR2 (N2858, N2857, N2630);
nand NAND4 (N2859, N2848, N1222, N922, N1475);
xor XOR2 (N2860, N2850, N2467);
nor NOR2 (N2861, N2855, N255);
or OR2 (N2862, N2856, N977);
or OR3 (N2863, N2854, N840, N943);
nand NAND4 (N2864, N2846, N907, N1378, N665);
nor NOR3 (N2865, N2849, N61, N883);
xor XOR2 (N2866, N2858, N1077);
not NOT1 (N2867, N2865);
nand NAND2 (N2868, N2867, N1596);
nor NOR2 (N2869, N2845, N1236);
nor NOR3 (N2870, N2868, N2659, N1526);
nand NAND4 (N2871, N2863, N809, N244, N2270);
nor NOR3 (N2872, N2864, N657, N904);
nand NAND3 (N2873, N2866, N932, N672);
nor NOR3 (N2874, N2869, N1553, N2422);
not NOT1 (N2875, N2870);
and AND4 (N2876, N2860, N2700, N299, N1658);
xor XOR2 (N2877, N2871, N1322);
and AND4 (N2878, N2876, N2086, N1059, N1751);
and AND2 (N2879, N2859, N2399);
and AND3 (N2880, N2862, N2838, N1220);
not NOT1 (N2881, N2880);
and AND3 (N2882, N2873, N2849, N1285);
or OR2 (N2883, N2852, N1682);
buf BUF1 (N2884, N2882);
xor XOR2 (N2885, N2878, N1569);
and AND3 (N2886, N2874, N2234, N1062);
or OR2 (N2887, N2881, N915);
nand NAND4 (N2888, N2872, N630, N393, N2084);
and AND4 (N2889, N2861, N156, N2091, N2721);
and AND4 (N2890, N2888, N615, N1590, N2566);
xor XOR2 (N2891, N2885, N564);
buf BUF1 (N2892, N2887);
not NOT1 (N2893, N2889);
buf BUF1 (N2894, N2877);
xor XOR2 (N2895, N2884, N2628);
or OR4 (N2896, N2886, N1928, N2816, N164);
or OR4 (N2897, N2896, N2162, N1084, N1769);
and AND3 (N2898, N2875, N1688, N1792);
nor NOR3 (N2899, N2894, N1470, N902);
and AND4 (N2900, N2898, N696, N115, N417);
or OR2 (N2901, N2890, N1231);
and AND2 (N2902, N2901, N511);
nor NOR3 (N2903, N2891, N2690, N517);
and AND4 (N2904, N2902, N2227, N1952, N1992);
buf BUF1 (N2905, N2893);
and AND3 (N2906, N2903, N2727, N1629);
and AND3 (N2907, N2906, N2305, N1882);
not NOT1 (N2908, N2907);
nor NOR3 (N2909, N2895, N1267, N2642);
nand NAND3 (N2910, N2908, N2424, N1121);
or OR4 (N2911, N2879, N2193, N2460, N557);
and AND2 (N2912, N2904, N2283);
xor XOR2 (N2913, N2912, N1434);
nand NAND3 (N2914, N2905, N801, N1463);
nand NAND4 (N2915, N2911, N442, N1167, N2059);
xor XOR2 (N2916, N2915, N2177);
nor NOR3 (N2917, N2914, N2643, N1308);
xor XOR2 (N2918, N2917, N2886);
xor XOR2 (N2919, N2909, N2405);
or OR3 (N2920, N2899, N1595, N1684);
buf BUF1 (N2921, N2892);
or OR2 (N2922, N2897, N115);
and AND2 (N2923, N2918, N1472);
and AND3 (N2924, N2910, N2320, N198);
or OR2 (N2925, N2921, N1837);
xor XOR2 (N2926, N2883, N731);
xor XOR2 (N2927, N2925, N535);
and AND2 (N2928, N2924, N1317);
and AND3 (N2929, N2916, N2666, N1856);
nand NAND3 (N2930, N2919, N1781, N736);
buf BUF1 (N2931, N2920);
or OR4 (N2932, N2931, N1908, N1330, N2276);
or OR3 (N2933, N2900, N70, N1720);
and AND2 (N2934, N2927, N2816);
nand NAND3 (N2935, N2913, N1773, N1806);
xor XOR2 (N2936, N2935, N1665);
xor XOR2 (N2937, N2930, N2000);
and AND2 (N2938, N2936, N2578);
and AND4 (N2939, N2929, N2845, N2222, N1045);
xor XOR2 (N2940, N2938, N1909);
and AND2 (N2941, N2928, N570);
not NOT1 (N2942, N2932);
not NOT1 (N2943, N2933);
buf BUF1 (N2944, N2934);
xor XOR2 (N2945, N2942, N28);
buf BUF1 (N2946, N2943);
nor NOR3 (N2947, N2937, N2491, N109);
nor NOR2 (N2948, N2941, N522);
and AND3 (N2949, N2940, N1545, N1744);
buf BUF1 (N2950, N2926);
and AND4 (N2951, N2947, N293, N2411, N524);
nand NAND4 (N2952, N2946, N2357, N2639, N2599);
nor NOR3 (N2953, N2948, N1959, N1055);
buf BUF1 (N2954, N2923);
nand NAND2 (N2955, N2953, N592);
buf BUF1 (N2956, N2954);
or OR3 (N2957, N2922, N431, N948);
xor XOR2 (N2958, N2955, N2697);
nand NAND2 (N2959, N2956, N2427);
buf BUF1 (N2960, N2939);
or OR2 (N2961, N2952, N2408);
buf BUF1 (N2962, N2950);
xor XOR2 (N2963, N2960, N1034);
and AND3 (N2964, N2945, N1523, N2758);
not NOT1 (N2965, N2951);
buf BUF1 (N2966, N2964);
nand NAND3 (N2967, N2957, N392, N1277);
not NOT1 (N2968, N2959);
nor NOR4 (N2969, N2963, N646, N2069, N2328);
and AND3 (N2970, N2961, N496, N2280);
not NOT1 (N2971, N2949);
buf BUF1 (N2972, N2962);
and AND4 (N2973, N2969, N2942, N626, N2138);
and AND4 (N2974, N2968, N174, N824, N1231);
nor NOR3 (N2975, N2970, N506, N2956);
xor XOR2 (N2976, N2973, N1203);
or OR3 (N2977, N2971, N1689, N535);
nand NAND2 (N2978, N2965, N1681);
buf BUF1 (N2979, N2974);
or OR2 (N2980, N2966, N2403);
buf BUF1 (N2981, N2967);
and AND3 (N2982, N2977, N1004, N2531);
nand NAND2 (N2983, N2979, N651);
or OR4 (N2984, N2944, N61, N121, N2946);
or OR2 (N2985, N2982, N40);
not NOT1 (N2986, N2980);
buf BUF1 (N2987, N2981);
not NOT1 (N2988, N2987);
not NOT1 (N2989, N2958);
buf BUF1 (N2990, N2972);
and AND2 (N2991, N2978, N1997);
or OR3 (N2992, N2991, N2968, N2027);
buf BUF1 (N2993, N2990);
or OR2 (N2994, N2975, N1694);
or OR3 (N2995, N2985, N2521, N1760);
xor XOR2 (N2996, N2989, N1663);
nand NAND3 (N2997, N2996, N1227, N2201);
nand NAND2 (N2998, N2993, N1061);
not NOT1 (N2999, N2988);
not NOT1 (N3000, N2999);
nand NAND4 (N3001, N2992, N2471, N639, N2966);
buf BUF1 (N3002, N2995);
and AND2 (N3003, N2976, N1028);
buf BUF1 (N3004, N2998);
nor NOR3 (N3005, N3001, N840, N184);
not NOT1 (N3006, N3005);
nand NAND4 (N3007, N3004, N520, N329, N218);
not NOT1 (N3008, N2986);
or OR4 (N3009, N3003, N2781, N652, N1277);
or OR4 (N3010, N3000, N1785, N523, N478);
nand NAND2 (N3011, N3002, N1918);
and AND3 (N3012, N3010, N1336, N2779);
nand NAND4 (N3013, N3011, N1133, N1782, N2350);
nand NAND2 (N3014, N3008, N2469);
xor XOR2 (N3015, N3012, N1652);
buf BUF1 (N3016, N2994);
and AND3 (N3017, N2983, N2353, N3001);
and AND4 (N3018, N2997, N2424, N1002, N2978);
or OR4 (N3019, N3013, N1978, N1008, N1176);
nand NAND2 (N3020, N3018, N1080);
xor XOR2 (N3021, N3007, N505);
or OR2 (N3022, N3006, N1077);
nor NOR2 (N3023, N3019, N99);
nor NOR3 (N3024, N3021, N856, N1791);
xor XOR2 (N3025, N3023, N179);
nand NAND3 (N3026, N3014, N389, N2416);
not NOT1 (N3027, N3026);
not NOT1 (N3028, N3017);
or OR3 (N3029, N3016, N2733, N1214);
and AND3 (N3030, N3024, N679, N780);
nand NAND3 (N3031, N3030, N48, N1466);
nand NAND3 (N3032, N3028, N124, N94);
and AND2 (N3033, N3020, N2425);
or OR2 (N3034, N3009, N1881);
and AND2 (N3035, N3029, N2550);
xor XOR2 (N3036, N3035, N466);
nand NAND3 (N3037, N3022, N2108, N2821);
xor XOR2 (N3038, N3027, N2414);
nand NAND4 (N3039, N3036, N1414, N2936, N2985);
nand NAND3 (N3040, N3038, N1612, N162);
or OR4 (N3041, N3039, N2703, N192, N2897);
xor XOR2 (N3042, N3015, N3015);
and AND4 (N3043, N3033, N2770, N1424, N994);
nor NOR3 (N3044, N2984, N862, N1912);
and AND2 (N3045, N3044, N2698);
or OR4 (N3046, N3041, N1803, N493, N2801);
xor XOR2 (N3047, N3037, N2052);
nand NAND2 (N3048, N3031, N862);
not NOT1 (N3049, N3043);
and AND2 (N3050, N3048, N433);
nand NAND4 (N3051, N3046, N899, N260, N1072);
buf BUF1 (N3052, N3034);
nand NAND4 (N3053, N3025, N439, N596, N2415);
nand NAND4 (N3054, N3050, N334, N1864, N1033);
or OR2 (N3055, N3053, N715);
and AND4 (N3056, N3055, N2392, N2117, N2641);
nor NOR4 (N3057, N3042, N2779, N2234, N2976);
buf BUF1 (N3058, N3049);
xor XOR2 (N3059, N3051, N1577);
nand NAND4 (N3060, N3057, N2100, N2828, N1798);
nand NAND3 (N3061, N3060, N2891, N2847);
or OR3 (N3062, N3061, N1767, N260);
or OR2 (N3063, N3056, N1065);
nor NOR4 (N3064, N3047, N1708, N1342, N554);
not NOT1 (N3065, N3045);
nand NAND4 (N3066, N3059, N927, N300, N2340);
xor XOR2 (N3067, N3063, N1812);
xor XOR2 (N3068, N3066, N2696);
or OR3 (N3069, N3052, N983, N582);
nand NAND4 (N3070, N3058, N2781, N163, N1767);
buf BUF1 (N3071, N3065);
and AND4 (N3072, N3069, N1112, N2683, N2155);
nand NAND4 (N3073, N3040, N1198, N1517, N1334);
buf BUF1 (N3074, N3054);
nand NAND3 (N3075, N3074, N62, N2413);
nand NAND2 (N3076, N3071, N192);
nor NOR4 (N3077, N3068, N2244, N1104, N1649);
not NOT1 (N3078, N3077);
and AND2 (N3079, N3062, N1288);
nand NAND3 (N3080, N3075, N2057, N1754);
nand NAND4 (N3081, N3067, N3045, N1450, N2234);
nand NAND4 (N3082, N3076, N1188, N3002, N2106);
and AND4 (N3083, N3072, N699, N1125, N998);
and AND4 (N3084, N3079, N2976, N902, N1250);
xor XOR2 (N3085, N3078, N894);
or OR2 (N3086, N3083, N2318);
not NOT1 (N3087, N3070);
not NOT1 (N3088, N3082);
buf BUF1 (N3089, N3073);
nand NAND2 (N3090, N3081, N187);
and AND3 (N3091, N3088, N2886, N2991);
buf BUF1 (N3092, N3091);
nand NAND2 (N3093, N3032, N1388);
not NOT1 (N3094, N3064);
nand NAND2 (N3095, N3086, N1662);
or OR2 (N3096, N3095, N578);
nand NAND3 (N3097, N3084, N2151, N1145);
xor XOR2 (N3098, N3085, N798);
not NOT1 (N3099, N3094);
nand NAND4 (N3100, N3089, N503, N1989, N2303);
nor NOR2 (N3101, N3100, N143);
or OR4 (N3102, N3101, N1930, N2519, N2994);
nand NAND3 (N3103, N3102, N1012, N44);
nor NOR4 (N3104, N3087, N551, N2185, N1794);
and AND2 (N3105, N3096, N683);
and AND4 (N3106, N3103, N678, N1978, N2704);
nor NOR2 (N3107, N3106, N41);
nor NOR3 (N3108, N3104, N2710, N1736);
nor NOR3 (N3109, N3097, N1363, N2031);
or OR3 (N3110, N3107, N1918, N2772);
buf BUF1 (N3111, N3108);
and AND4 (N3112, N3090, N722, N1315, N2574);
buf BUF1 (N3113, N3099);
not NOT1 (N3114, N3092);
or OR3 (N3115, N3080, N2216, N1443);
or OR4 (N3116, N3111, N2186, N2593, N872);
xor XOR2 (N3117, N3109, N596);
xor XOR2 (N3118, N3113, N1775);
buf BUF1 (N3119, N3115);
nand NAND2 (N3120, N3114, N374);
buf BUF1 (N3121, N3119);
nor NOR3 (N3122, N3117, N2262, N1643);
or OR3 (N3123, N3121, N216, N1999);
not NOT1 (N3124, N3110);
buf BUF1 (N3125, N3122);
buf BUF1 (N3126, N3116);
xor XOR2 (N3127, N3093, N2640);
nand NAND4 (N3128, N3123, N536, N2521, N3017);
and AND3 (N3129, N3098, N2949, N1257);
buf BUF1 (N3130, N3128);
and AND4 (N3131, N3126, N1164, N2091, N663);
nor NOR4 (N3132, N3120, N2493, N2581, N1299);
nand NAND3 (N3133, N3105, N2303, N2947);
xor XOR2 (N3134, N3133, N2560);
and AND4 (N3135, N3129, N1025, N36, N1265);
xor XOR2 (N3136, N3132, N1706);
and AND2 (N3137, N3127, N1145);
nand NAND2 (N3138, N3135, N649);
and AND2 (N3139, N3131, N2444);
or OR2 (N3140, N3118, N2360);
buf BUF1 (N3141, N3125);
not NOT1 (N3142, N3140);
nor NOR3 (N3143, N3124, N2475, N1220);
or OR2 (N3144, N3138, N2226);
nor NOR4 (N3145, N3112, N771, N2117, N2596);
xor XOR2 (N3146, N3142, N1600);
xor XOR2 (N3147, N3143, N2663);
nand NAND4 (N3148, N3130, N789, N3019, N140);
buf BUF1 (N3149, N3141);
buf BUF1 (N3150, N3144);
buf BUF1 (N3151, N3139);
buf BUF1 (N3152, N3145);
nand NAND2 (N3153, N3152, N712);
and AND3 (N3154, N3149, N991, N2084);
xor XOR2 (N3155, N3148, N133);
nand NAND2 (N3156, N3136, N1519);
and AND4 (N3157, N3155, N2526, N1497, N1156);
or OR2 (N3158, N3147, N1647);
not NOT1 (N3159, N3157);
xor XOR2 (N3160, N3137, N3071);
not NOT1 (N3161, N3156);
nor NOR2 (N3162, N3134, N1653);
not NOT1 (N3163, N3151);
not NOT1 (N3164, N3160);
not NOT1 (N3165, N3161);
or OR3 (N3166, N3159, N1279, N1792);
and AND2 (N3167, N3150, N2792);
nor NOR3 (N3168, N3164, N682, N2838);
nand NAND4 (N3169, N3163, N1882, N2108, N2526);
not NOT1 (N3170, N3169);
not NOT1 (N3171, N3146);
not NOT1 (N3172, N3153);
and AND4 (N3173, N3167, N1944, N1379, N1485);
xor XOR2 (N3174, N3158, N1315);
buf BUF1 (N3175, N3172);
not NOT1 (N3176, N3170);
nor NOR3 (N3177, N3165, N2399, N373);
nor NOR2 (N3178, N3174, N1462);
nor NOR4 (N3179, N3178, N1791, N2549, N2845);
xor XOR2 (N3180, N3171, N19);
nor NOR2 (N3181, N3175, N777);
xor XOR2 (N3182, N3177, N70);
and AND3 (N3183, N3168, N1270, N790);
nor NOR4 (N3184, N3173, N1747, N1086, N1374);
buf BUF1 (N3185, N3180);
buf BUF1 (N3186, N3183);
not NOT1 (N3187, N3154);
and AND3 (N3188, N3181, N2639, N2093);
nor NOR2 (N3189, N3162, N1984);
xor XOR2 (N3190, N3176, N188);
not NOT1 (N3191, N3186);
not NOT1 (N3192, N3191);
not NOT1 (N3193, N3179);
xor XOR2 (N3194, N3187, N2215);
nor NOR2 (N3195, N3185, N2218);
buf BUF1 (N3196, N3182);
xor XOR2 (N3197, N3195, N1955);
nand NAND3 (N3198, N3193, N405, N2739);
buf BUF1 (N3199, N3190);
nand NAND3 (N3200, N3198, N2435, N1671);
nand NAND3 (N3201, N3200, N95, N720);
nor NOR2 (N3202, N3199, N3092);
or OR4 (N3203, N3201, N2751, N2646, N2740);
buf BUF1 (N3204, N3203);
xor XOR2 (N3205, N3192, N2181);
buf BUF1 (N3206, N3202);
not NOT1 (N3207, N3189);
xor XOR2 (N3208, N3166, N1888);
nand NAND4 (N3209, N3208, N2806, N364, N2334);
nand NAND4 (N3210, N3204, N1212, N45, N132);
buf BUF1 (N3211, N3184);
nand NAND2 (N3212, N3194, N761);
and AND2 (N3213, N3205, N2927);
buf BUF1 (N3214, N3207);
and AND2 (N3215, N3206, N2915);
or OR2 (N3216, N3211, N2720);
or OR3 (N3217, N3188, N860, N3036);
nor NOR2 (N3218, N3217, N386);
and AND2 (N3219, N3209, N30);
buf BUF1 (N3220, N3213);
xor XOR2 (N3221, N3214, N3120);
nor NOR4 (N3222, N3215, N1608, N2365, N292);
xor XOR2 (N3223, N3218, N3041);
and AND3 (N3224, N3221, N5, N1822);
not NOT1 (N3225, N3224);
nor NOR4 (N3226, N3223, N2500, N2140, N300);
and AND4 (N3227, N3212, N2991, N554, N2132);
buf BUF1 (N3228, N3210);
and AND3 (N3229, N3226, N2241, N496);
and AND3 (N3230, N3228, N437, N575);
xor XOR2 (N3231, N3230, N374);
or OR2 (N3232, N3225, N1768);
nor NOR2 (N3233, N3196, N935);
or OR4 (N3234, N3220, N2992, N1493, N1606);
not NOT1 (N3235, N3222);
and AND3 (N3236, N3231, N209, N1264);
buf BUF1 (N3237, N3235);
and AND4 (N3238, N3236, N1356, N1524, N2077);
not NOT1 (N3239, N3229);
not NOT1 (N3240, N3234);
and AND2 (N3241, N3232, N135);
and AND3 (N3242, N3241, N2648, N2822);
and AND4 (N3243, N3237, N1588, N3007, N471);
nor NOR3 (N3244, N3240, N2350, N1901);
and AND3 (N3245, N3227, N816, N275);
and AND4 (N3246, N3197, N2585, N139, N908);
buf BUF1 (N3247, N3246);
xor XOR2 (N3248, N3247, N874);
xor XOR2 (N3249, N3248, N1244);
nand NAND3 (N3250, N3219, N1101, N1550);
nand NAND2 (N3251, N3238, N259);
xor XOR2 (N3252, N3243, N2656);
and AND4 (N3253, N3252, N3074, N2906, N715);
and AND2 (N3254, N3253, N2625);
xor XOR2 (N3255, N3254, N1034);
not NOT1 (N3256, N3216);
nand NAND2 (N3257, N3245, N1139);
xor XOR2 (N3258, N3244, N2817);
or OR4 (N3259, N3239, N235, N868, N474);
nand NAND2 (N3260, N3259, N2266);
nand NAND2 (N3261, N3242, N1905);
not NOT1 (N3262, N3257);
buf BUF1 (N3263, N3233);
xor XOR2 (N3264, N3250, N243);
and AND4 (N3265, N3260, N1918, N1083, N2814);
buf BUF1 (N3266, N3255);
or OR2 (N3267, N3264, N1636);
or OR3 (N3268, N3251, N1216, N2911);
and AND4 (N3269, N3256, N2860, N1003, N2508);
nand NAND2 (N3270, N3269, N1593);
nand NAND4 (N3271, N3265, N2635, N129, N703);
not NOT1 (N3272, N3249);
buf BUF1 (N3273, N3266);
buf BUF1 (N3274, N3263);
buf BUF1 (N3275, N3270);
nor NOR2 (N3276, N3273, N2465);
and AND4 (N3277, N3261, N922, N3199, N3271);
nor NOR3 (N3278, N381, N2790, N1538);
nor NOR3 (N3279, N3276, N1924, N132);
nand NAND3 (N3280, N3272, N2346, N2249);
buf BUF1 (N3281, N3279);
or OR2 (N3282, N3278, N680);
buf BUF1 (N3283, N3258);
nor NOR3 (N3284, N3277, N750, N762);
and AND4 (N3285, N3282, N641, N1048, N2050);
nor NOR4 (N3286, N3285, N2290, N2989, N2510);
not NOT1 (N3287, N3281);
not NOT1 (N3288, N3286);
buf BUF1 (N3289, N3275);
buf BUF1 (N3290, N3289);
xor XOR2 (N3291, N3283, N1163);
nand NAND4 (N3292, N3280, N2919, N1034, N3172);
nand NAND3 (N3293, N3288, N1553, N1698);
not NOT1 (N3294, N3284);
nor NOR2 (N3295, N3274, N1076);
nand NAND3 (N3296, N3292, N512, N584);
nand NAND2 (N3297, N3294, N3088);
xor XOR2 (N3298, N3290, N2868);
nand NAND2 (N3299, N3293, N2490);
buf BUF1 (N3300, N3298);
and AND2 (N3301, N3299, N348);
nor NOR2 (N3302, N3295, N2191);
nor NOR3 (N3303, N3297, N154, N2369);
not NOT1 (N3304, N3301);
nand NAND3 (N3305, N3296, N1429, N89);
nand NAND4 (N3306, N3305, N2424, N2375, N2627);
nand NAND4 (N3307, N3306, N2567, N2712, N1132);
xor XOR2 (N3308, N3287, N3054);
nor NOR3 (N3309, N3300, N2936, N1833);
buf BUF1 (N3310, N3309);
xor XOR2 (N3311, N3291, N1648);
and AND3 (N3312, N3267, N571, N595);
and AND2 (N3313, N3308, N1268);
xor XOR2 (N3314, N3303, N496);
or OR3 (N3315, N3307, N256, N2421);
buf BUF1 (N3316, N3315);
and AND3 (N3317, N3316, N51, N1374);
nand NAND3 (N3318, N3317, N1383, N1390);
and AND4 (N3319, N3268, N2822, N1293, N540);
not NOT1 (N3320, N3302);
nor NOR3 (N3321, N3304, N263, N1789);
xor XOR2 (N3322, N3321, N1980);
nand NAND2 (N3323, N3314, N82);
or OR2 (N3324, N3320, N2297);
not NOT1 (N3325, N3324);
buf BUF1 (N3326, N3319);
and AND2 (N3327, N3310, N2956);
xor XOR2 (N3328, N3322, N1706);
nor NOR4 (N3329, N3313, N155, N2031, N755);
or OR3 (N3330, N3326, N2404, N413);
buf BUF1 (N3331, N3328);
nor NOR4 (N3332, N3327, N3185, N2811, N2033);
not NOT1 (N3333, N3323);
and AND4 (N3334, N3311, N2708, N999, N1829);
nor NOR3 (N3335, N3329, N3258, N1994);
not NOT1 (N3336, N3334);
nand NAND2 (N3337, N3312, N2762);
and AND3 (N3338, N3335, N416, N910);
xor XOR2 (N3339, N3262, N814);
and AND2 (N3340, N3337, N1879);
or OR2 (N3341, N3340, N2832);
and AND2 (N3342, N3318, N2392);
buf BUF1 (N3343, N3333);
and AND2 (N3344, N3331, N2192);
nand NAND2 (N3345, N3336, N2673);
xor XOR2 (N3346, N3345, N208);
nand NAND3 (N3347, N3332, N2186, N586);
and AND4 (N3348, N3346, N2867, N931, N737);
nand NAND2 (N3349, N3341, N757);
nor NOR2 (N3350, N3348, N2639);
and AND4 (N3351, N3330, N1624, N2725, N2845);
not NOT1 (N3352, N3344);
nor NOR4 (N3353, N3342, N2038, N903, N827);
nor NOR4 (N3354, N3353, N150, N3062, N1544);
nor NOR3 (N3355, N3339, N3210, N738);
not NOT1 (N3356, N3338);
xor XOR2 (N3357, N3349, N1078);
nor NOR4 (N3358, N3357, N891, N3168, N2553);
or OR3 (N3359, N3356, N3308, N1229);
or OR4 (N3360, N3343, N2577, N11, N3284);
buf BUF1 (N3361, N3354);
not NOT1 (N3362, N3350);
nor NOR2 (N3363, N3362, N2912);
and AND2 (N3364, N3351, N245);
or OR2 (N3365, N3359, N1360);
buf BUF1 (N3366, N3325);
nand NAND4 (N3367, N3352, N2279, N2684, N3142);
buf BUF1 (N3368, N3358);
buf BUF1 (N3369, N3360);
xor XOR2 (N3370, N3365, N2548);
or OR2 (N3371, N3364, N1571);
buf BUF1 (N3372, N3367);
nor NOR2 (N3373, N3372, N1295);
nor NOR3 (N3374, N3361, N27, N1811);
and AND4 (N3375, N3370, N1755, N20, N664);
or OR3 (N3376, N3374, N69, N585);
nand NAND2 (N3377, N3347, N3341);
or OR3 (N3378, N3373, N2814, N180);
and AND3 (N3379, N3378, N2768, N3271);
nand NAND2 (N3380, N3377, N2086);
buf BUF1 (N3381, N3376);
buf BUF1 (N3382, N3368);
nor NOR2 (N3383, N3369, N3270);
or OR4 (N3384, N3380, N798, N1166, N3201);
xor XOR2 (N3385, N3379, N882);
or OR3 (N3386, N3381, N1750, N1872);
and AND3 (N3387, N3383, N2592, N2671);
buf BUF1 (N3388, N3366);
xor XOR2 (N3389, N3385, N3353);
nor NOR3 (N3390, N3355, N1769, N1573);
nand NAND2 (N3391, N3371, N2053);
xor XOR2 (N3392, N3390, N2920);
not NOT1 (N3393, N3363);
buf BUF1 (N3394, N3393);
not NOT1 (N3395, N3388);
nor NOR2 (N3396, N3386, N2769);
not NOT1 (N3397, N3394);
not NOT1 (N3398, N3375);
not NOT1 (N3399, N3398);
nor NOR3 (N3400, N3397, N2082, N2755);
nand NAND2 (N3401, N3382, N1978);
not NOT1 (N3402, N3401);
buf BUF1 (N3403, N3387);
nand NAND2 (N3404, N3392, N469);
xor XOR2 (N3405, N3402, N3136);
buf BUF1 (N3406, N3389);
nand NAND3 (N3407, N3406, N1569, N3227);
and AND2 (N3408, N3384, N36);
and AND4 (N3409, N3395, N1949, N3186, N1075);
nand NAND3 (N3410, N3396, N885, N2154);
xor XOR2 (N3411, N3410, N2155);
and AND3 (N3412, N3408, N1200, N2579);
nand NAND3 (N3413, N3399, N2932, N815);
not NOT1 (N3414, N3400);
xor XOR2 (N3415, N3391, N1869);
nor NOR3 (N3416, N3405, N2508, N3188);
xor XOR2 (N3417, N3416, N2005);
nand NAND3 (N3418, N3412, N748, N185);
or OR4 (N3419, N3404, N2250, N1473, N3289);
nand NAND4 (N3420, N3415, N2896, N1454, N3213);
buf BUF1 (N3421, N3413);
and AND4 (N3422, N3417, N2234, N1820, N388);
not NOT1 (N3423, N3409);
buf BUF1 (N3424, N3423);
or OR4 (N3425, N3422, N2214, N2937, N2281);
not NOT1 (N3426, N3403);
or OR4 (N3427, N3424, N2464, N831, N495);
nand NAND3 (N3428, N3418, N2814, N3012);
nor NOR4 (N3429, N3407, N1295, N2822, N3314);
and AND3 (N3430, N3428, N907, N1758);
or OR3 (N3431, N3414, N1079, N2011);
nor NOR4 (N3432, N3431, N598, N2987, N478);
or OR4 (N3433, N3432, N1833, N1428, N1274);
not NOT1 (N3434, N3419);
nor NOR2 (N3435, N3425, N1974);
nand NAND4 (N3436, N3421, N2614, N735, N3039);
nor NOR4 (N3437, N3420, N2224, N1773, N1282);
nand NAND3 (N3438, N3436, N1873, N684);
not NOT1 (N3439, N3430);
nand NAND4 (N3440, N3433, N295, N2610, N2359);
not NOT1 (N3441, N3426);
and AND4 (N3442, N3439, N2438, N1774, N1149);
not NOT1 (N3443, N3429);
nand NAND4 (N3444, N3441, N872, N1378, N1341);
xor XOR2 (N3445, N3434, N1759);
nand NAND3 (N3446, N3444, N441, N31);
xor XOR2 (N3447, N3437, N1553);
xor XOR2 (N3448, N3446, N3276);
xor XOR2 (N3449, N3445, N1568);
not NOT1 (N3450, N3438);
or OR3 (N3451, N3440, N3334, N1521);
or OR2 (N3452, N3427, N449);
xor XOR2 (N3453, N3450, N783);
xor XOR2 (N3454, N3453, N696);
nand NAND4 (N3455, N3448, N1586, N2214, N526);
xor XOR2 (N3456, N3454, N1182);
xor XOR2 (N3457, N3449, N2581);
nor NOR4 (N3458, N3443, N3216, N2167, N3030);
nand NAND3 (N3459, N3435, N303, N3211);
xor XOR2 (N3460, N3447, N668);
nand NAND2 (N3461, N3455, N3207);
nand NAND2 (N3462, N3451, N2300);
xor XOR2 (N3463, N3459, N435);
not NOT1 (N3464, N3457);
or OR4 (N3465, N3461, N3309, N966, N504);
nor NOR2 (N3466, N3464, N3005);
nor NOR4 (N3467, N3456, N3262, N784, N1396);
or OR3 (N3468, N3452, N3389, N716);
and AND2 (N3469, N3460, N752);
and AND4 (N3470, N3469, N997, N1616, N610);
buf BUF1 (N3471, N3442);
xor XOR2 (N3472, N3458, N199);
nand NAND3 (N3473, N3462, N872, N997);
and AND4 (N3474, N3472, N3373, N2664, N150);
buf BUF1 (N3475, N3467);
nand NAND2 (N3476, N3471, N1348);
xor XOR2 (N3477, N3473, N802);
nor NOR4 (N3478, N3474, N2760, N2271, N2378);
buf BUF1 (N3479, N3465);
buf BUF1 (N3480, N3466);
or OR4 (N3481, N3411, N1608, N7, N1385);
xor XOR2 (N3482, N3478, N908);
not NOT1 (N3483, N3476);
and AND3 (N3484, N3480, N1050, N51);
buf BUF1 (N3485, N3481);
xor XOR2 (N3486, N3482, N2667);
nor NOR4 (N3487, N3477, N1987, N3461, N3385);
and AND3 (N3488, N3470, N1828, N3162);
and AND2 (N3489, N3484, N327);
xor XOR2 (N3490, N3479, N363);
xor XOR2 (N3491, N3486, N66);
nand NAND3 (N3492, N3491, N1180, N2037);
xor XOR2 (N3493, N3463, N2202);
buf BUF1 (N3494, N3490);
nor NOR4 (N3495, N3485, N1383, N2358, N1817);
nor NOR2 (N3496, N3495, N1076);
xor XOR2 (N3497, N3494, N602);
nor NOR2 (N3498, N3483, N2643);
nor NOR3 (N3499, N3493, N587, N361);
or OR4 (N3500, N3468, N2233, N694, N1682);
nand NAND3 (N3501, N3475, N2452, N2062);
nor NOR4 (N3502, N3492, N2940, N2865, N1389);
or OR4 (N3503, N3488, N1281, N2676, N1269);
not NOT1 (N3504, N3489);
or OR2 (N3505, N3487, N2643);
buf BUF1 (N3506, N3500);
nor NOR4 (N3507, N3503, N212, N676, N269);
and AND2 (N3508, N3496, N2567);
and AND3 (N3509, N3497, N869, N531);
and AND3 (N3510, N3501, N2689, N328);
not NOT1 (N3511, N3504);
buf BUF1 (N3512, N3507);
not NOT1 (N3513, N3509);
xor XOR2 (N3514, N3511, N3409);
not NOT1 (N3515, N3505);
not NOT1 (N3516, N3515);
not NOT1 (N3517, N3499);
and AND2 (N3518, N3516, N2628);
not NOT1 (N3519, N3513);
not NOT1 (N3520, N3517);
or OR4 (N3521, N3510, N807, N66, N1597);
buf BUF1 (N3522, N3502);
not NOT1 (N3523, N3498);
xor XOR2 (N3524, N3506, N2020);
or OR2 (N3525, N3520, N940);
nand NAND3 (N3526, N3508, N3522, N478);
nand NAND3 (N3527, N3040, N2153, N3297);
xor XOR2 (N3528, N3527, N2608);
nor NOR3 (N3529, N3523, N2909, N2234);
or OR4 (N3530, N3525, N3337, N2275, N1037);
not NOT1 (N3531, N3512);
nand NAND2 (N3532, N3526, N44);
nand NAND3 (N3533, N3531, N2894, N1213);
nor NOR3 (N3534, N3518, N299, N3009);
and AND3 (N3535, N3533, N2819, N1304);
and AND2 (N3536, N3528, N2508);
nor NOR3 (N3537, N3519, N1661, N591);
not NOT1 (N3538, N3532);
buf BUF1 (N3539, N3537);
not NOT1 (N3540, N3530);
and AND2 (N3541, N3535, N2043);
xor XOR2 (N3542, N3539, N2704);
buf BUF1 (N3543, N3529);
nand NAND4 (N3544, N3541, N2267, N119, N1064);
xor XOR2 (N3545, N3538, N3426);
or OR2 (N3546, N3534, N2088);
buf BUF1 (N3547, N3542);
nand NAND3 (N3548, N3524, N11, N1150);
buf BUF1 (N3549, N3540);
nor NOR4 (N3550, N3521, N2299, N3525, N888);
buf BUF1 (N3551, N3548);
or OR2 (N3552, N3550, N1691);
and AND4 (N3553, N3544, N1154, N1066, N628);
xor XOR2 (N3554, N3546, N2837);
or OR2 (N3555, N3549, N2990);
xor XOR2 (N3556, N3555, N1024);
not NOT1 (N3557, N3554);
xor XOR2 (N3558, N3553, N754);
and AND2 (N3559, N3543, N2347);
nor NOR2 (N3560, N3559, N122);
nand NAND3 (N3561, N3552, N92, N1613);
and AND4 (N3562, N3557, N20, N47, N1392);
buf BUF1 (N3563, N3562);
xor XOR2 (N3564, N3545, N2331);
nor NOR3 (N3565, N3558, N693, N1898);
xor XOR2 (N3566, N3514, N1174);
not NOT1 (N3567, N3565);
not NOT1 (N3568, N3564);
or OR4 (N3569, N3560, N3204, N3345, N1754);
xor XOR2 (N3570, N3568, N1868);
not NOT1 (N3571, N3551);
xor XOR2 (N3572, N3570, N465);
and AND4 (N3573, N3567, N971, N1955, N27);
buf BUF1 (N3574, N3569);
nor NOR3 (N3575, N3563, N2855, N2303);
or OR4 (N3576, N3575, N2086, N1305, N1712);
or OR4 (N3577, N3547, N769, N152, N3087);
or OR2 (N3578, N3536, N811);
not NOT1 (N3579, N3577);
or OR3 (N3580, N3561, N2883, N1917);
buf BUF1 (N3581, N3576);
nand NAND2 (N3582, N3579, N734);
and AND2 (N3583, N3581, N3052);
nor NOR2 (N3584, N3556, N2128);
or OR3 (N3585, N3584, N874, N391);
xor XOR2 (N3586, N3578, N121);
nand NAND4 (N3587, N3571, N433, N697, N720);
or OR3 (N3588, N3585, N2494, N1097);
xor XOR2 (N3589, N3587, N3111);
buf BUF1 (N3590, N3586);
not NOT1 (N3591, N3590);
nor NOR2 (N3592, N3574, N271);
xor XOR2 (N3593, N3580, N2406);
nor NOR2 (N3594, N3591, N1340);
not NOT1 (N3595, N3593);
nor NOR2 (N3596, N3595, N1180);
not NOT1 (N3597, N3588);
or OR2 (N3598, N3573, N3064);
nand NAND4 (N3599, N3592, N3433, N3210, N1496);
or OR3 (N3600, N3598, N1608, N417);
xor XOR2 (N3601, N3582, N1757);
nand NAND2 (N3602, N3566, N2316);
buf BUF1 (N3603, N3589);
or OR3 (N3604, N3600, N1404, N2024);
nand NAND2 (N3605, N3597, N2692);
buf BUF1 (N3606, N3596);
buf BUF1 (N3607, N3603);
buf BUF1 (N3608, N3594);
or OR2 (N3609, N3605, N163);
nand NAND2 (N3610, N3604, N2162);
and AND3 (N3611, N3610, N1815, N1062);
xor XOR2 (N3612, N3608, N915);
or OR2 (N3613, N3609, N2788);
xor XOR2 (N3614, N3572, N976);
not NOT1 (N3615, N3601);
buf BUF1 (N3616, N3611);
nand NAND4 (N3617, N3599, N2815, N335, N962);
buf BUF1 (N3618, N3616);
nand NAND4 (N3619, N3583, N2582, N2495, N2362);
and AND2 (N3620, N3612, N1180);
and AND2 (N3621, N3620, N13);
or OR4 (N3622, N3621, N2192, N1242, N603);
not NOT1 (N3623, N3618);
or OR2 (N3624, N3613, N660);
nand NAND3 (N3625, N3619, N1086, N1690);
and AND2 (N3626, N3615, N1369);
or OR2 (N3627, N3602, N2763);
not NOT1 (N3628, N3617);
buf BUF1 (N3629, N3623);
and AND2 (N3630, N3628, N1486);
nor NOR3 (N3631, N3624, N2486, N1341);
nor NOR4 (N3632, N3614, N1141, N495, N1552);
buf BUF1 (N3633, N3626);
xor XOR2 (N3634, N3622, N3354);
buf BUF1 (N3635, N3625);
and AND4 (N3636, N3629, N662, N2948, N501);
xor XOR2 (N3637, N3632, N655);
xor XOR2 (N3638, N3634, N158);
and AND4 (N3639, N3635, N3497, N1833, N1958);
buf BUF1 (N3640, N3638);
buf BUF1 (N3641, N3631);
nand NAND2 (N3642, N3640, N2739);
buf BUF1 (N3643, N3637);
or OR3 (N3644, N3636, N2323, N2249);
xor XOR2 (N3645, N3630, N556);
nand NAND3 (N3646, N3607, N3113, N36);
not NOT1 (N3647, N3645);
nand NAND3 (N3648, N3644, N3601, N379);
xor XOR2 (N3649, N3646, N332);
xor XOR2 (N3650, N3641, N2460);
nand NAND2 (N3651, N3642, N27);
not NOT1 (N3652, N3650);
and AND4 (N3653, N3606, N1442, N1077, N3548);
and AND4 (N3654, N3639, N3071, N2359, N2624);
nor NOR3 (N3655, N3653, N2392, N790);
xor XOR2 (N3656, N3633, N420);
and AND2 (N3657, N3643, N2657);
xor XOR2 (N3658, N3655, N2593);
and AND2 (N3659, N3648, N3336);
nor NOR2 (N3660, N3657, N2888);
not NOT1 (N3661, N3656);
not NOT1 (N3662, N3647);
and AND3 (N3663, N3627, N3488, N2610);
nor NOR4 (N3664, N3649, N514, N1663, N3498);
and AND4 (N3665, N3651, N2426, N2701, N3395);
xor XOR2 (N3666, N3665, N599);
nand NAND2 (N3667, N3664, N2423);
nand NAND4 (N3668, N3658, N848, N667, N3235);
not NOT1 (N3669, N3663);
nand NAND2 (N3670, N3669, N3387);
xor XOR2 (N3671, N3670, N2554);
nor NOR2 (N3672, N3660, N2265);
buf BUF1 (N3673, N3667);
buf BUF1 (N3674, N3654);
xor XOR2 (N3675, N3666, N300);
buf BUF1 (N3676, N3652);
nand NAND4 (N3677, N3676, N2060, N283, N1252);
nand NAND3 (N3678, N3673, N878, N2964);
buf BUF1 (N3679, N3662);
nor NOR4 (N3680, N3661, N3155, N2634, N1738);
and AND3 (N3681, N3679, N1888, N2548);
xor XOR2 (N3682, N3681, N815);
xor XOR2 (N3683, N3671, N1696);
buf BUF1 (N3684, N3674);
and AND4 (N3685, N3678, N1512, N1262, N2252);
and AND2 (N3686, N3677, N268);
xor XOR2 (N3687, N3680, N2915);
and AND4 (N3688, N3672, N2377, N892, N2440);
nor NOR2 (N3689, N3685, N2731);
or OR4 (N3690, N3659, N2286, N2447, N2490);
not NOT1 (N3691, N3690);
nor NOR3 (N3692, N3688, N3609, N1991);
not NOT1 (N3693, N3689);
nor NOR2 (N3694, N3693, N2615);
nor NOR2 (N3695, N3692, N2797);
nand NAND4 (N3696, N3683, N1557, N1268, N3278);
or OR4 (N3697, N3695, N601, N1262, N1639);
buf BUF1 (N3698, N3684);
not NOT1 (N3699, N3697);
and AND4 (N3700, N3696, N2549, N497, N1990);
and AND2 (N3701, N3687, N119);
nor NOR2 (N3702, N3668, N119);
nand NAND2 (N3703, N3699, N2191);
not NOT1 (N3704, N3675);
or OR4 (N3705, N3702, N61, N289, N327);
nand NAND4 (N3706, N3701, N2058, N2986, N3622);
xor XOR2 (N3707, N3704, N66);
or OR3 (N3708, N3706, N965, N2777);
not NOT1 (N3709, N3698);
nor NOR3 (N3710, N3682, N1889, N169);
and AND4 (N3711, N3705, N2227, N2042, N1166);
not NOT1 (N3712, N3710);
nand NAND4 (N3713, N3700, N615, N242, N487);
and AND3 (N3714, N3707, N3414, N681);
nand NAND4 (N3715, N3691, N1537, N1584, N738);
buf BUF1 (N3716, N3686);
nor NOR3 (N3717, N3712, N1139, N2999);
or OR3 (N3718, N3715, N431, N1844);
nand NAND2 (N3719, N3717, N2532);
and AND2 (N3720, N3709, N121);
or OR3 (N3721, N3713, N3717, N182);
nand NAND2 (N3722, N3708, N2872);
not NOT1 (N3723, N3716);
not NOT1 (N3724, N3719);
and AND2 (N3725, N3703, N1069);
not NOT1 (N3726, N3718);
or OR2 (N3727, N3725, N2528);
or OR3 (N3728, N3720, N1953, N3129);
not NOT1 (N3729, N3721);
buf BUF1 (N3730, N3694);
not NOT1 (N3731, N3730);
buf BUF1 (N3732, N3723);
xor XOR2 (N3733, N3731, N3550);
buf BUF1 (N3734, N3711);
buf BUF1 (N3735, N3734);
xor XOR2 (N3736, N3724, N240);
nand NAND3 (N3737, N3735, N807, N73);
or OR2 (N3738, N3726, N499);
nand NAND3 (N3739, N3733, N1948, N809);
not NOT1 (N3740, N3737);
buf BUF1 (N3741, N3727);
nand NAND3 (N3742, N3738, N924, N2428);
nand NAND3 (N3743, N3729, N3638, N621);
buf BUF1 (N3744, N3722);
not NOT1 (N3745, N3743);
and AND2 (N3746, N3741, N3336);
nand NAND4 (N3747, N3746, N2308, N2950, N282);
and AND4 (N3748, N3744, N1173, N1491, N3434);
not NOT1 (N3749, N3728);
nor NOR4 (N3750, N3749, N1891, N735, N1952);
and AND2 (N3751, N3732, N289);
xor XOR2 (N3752, N3747, N727);
nand NAND3 (N3753, N3748, N102, N100);
and AND3 (N3754, N3739, N2995, N2812);
or OR2 (N3755, N3742, N3210);
and AND2 (N3756, N3714, N3493);
nor NOR3 (N3757, N3750, N934, N1478);
or OR2 (N3758, N3751, N1430);
nand NAND2 (N3759, N3756, N1844);
nand NAND3 (N3760, N3759, N514, N112);
buf BUF1 (N3761, N3760);
nand NAND3 (N3762, N3745, N3049, N376);
not NOT1 (N3763, N3740);
nand NAND3 (N3764, N3755, N2883, N3280);
nor NOR2 (N3765, N3753, N1514);
buf BUF1 (N3766, N3763);
buf BUF1 (N3767, N3762);
or OR4 (N3768, N3764, N2588, N1457, N1696);
nand NAND2 (N3769, N3757, N2268);
not NOT1 (N3770, N3766);
xor XOR2 (N3771, N3765, N2486);
xor XOR2 (N3772, N3767, N132);
and AND4 (N3773, N3752, N3368, N73, N3275);
nand NAND2 (N3774, N3736, N958);
xor XOR2 (N3775, N3758, N1414);
xor XOR2 (N3776, N3768, N2206);
and AND4 (N3777, N3772, N1707, N2234, N2468);
or OR4 (N3778, N3773, N1565, N3616, N612);
or OR3 (N3779, N3774, N133, N883);
nor NOR3 (N3780, N3777, N2610, N834);
not NOT1 (N3781, N3761);
not NOT1 (N3782, N3779);
and AND2 (N3783, N3780, N3045);
not NOT1 (N3784, N3769);
nand NAND3 (N3785, N3770, N2848, N1179);
nor NOR4 (N3786, N3754, N1067, N2402, N202);
nor NOR3 (N3787, N3778, N1159, N2005);
xor XOR2 (N3788, N3782, N2840);
nor NOR4 (N3789, N3788, N2568, N738, N1611);
or OR2 (N3790, N3785, N719);
buf BUF1 (N3791, N3789);
xor XOR2 (N3792, N3787, N2156);
nand NAND3 (N3793, N3792, N3440, N99);
buf BUF1 (N3794, N3775);
buf BUF1 (N3795, N3781);
nand NAND4 (N3796, N3784, N3662, N693, N3285);
nor NOR2 (N3797, N3786, N1092);
buf BUF1 (N3798, N3791);
or OR3 (N3799, N3796, N177, N3189);
not NOT1 (N3800, N3771);
or OR3 (N3801, N3794, N607, N983);
buf BUF1 (N3802, N3783);
nor NOR3 (N3803, N3797, N571, N2338);
or OR2 (N3804, N3776, N419);
nand NAND4 (N3805, N3799, N3117, N1071, N1464);
or OR3 (N3806, N3805, N509, N311);
not NOT1 (N3807, N3800);
or OR4 (N3808, N3790, N3208, N1069, N1204);
nor NOR4 (N3809, N3806, N2088, N2126, N2237);
nor NOR2 (N3810, N3795, N2224);
nor NOR4 (N3811, N3804, N2569, N91, N779);
buf BUF1 (N3812, N3810);
or OR3 (N3813, N3793, N1149, N3711);
not NOT1 (N3814, N3807);
buf BUF1 (N3815, N3802);
not NOT1 (N3816, N3813);
buf BUF1 (N3817, N3814);
xor XOR2 (N3818, N3809, N3394);
nand NAND2 (N3819, N3816, N3650);
buf BUF1 (N3820, N3817);
nand NAND3 (N3821, N3808, N2747, N854);
buf BUF1 (N3822, N3818);
or OR2 (N3823, N3815, N1111);
xor XOR2 (N3824, N3812, N204);
xor XOR2 (N3825, N3819, N3002);
or OR2 (N3826, N3820, N1060);
nor NOR2 (N3827, N3801, N3315);
nand NAND4 (N3828, N3825, N1947, N3521, N384);
buf BUF1 (N3829, N3822);
and AND3 (N3830, N3798, N2844, N3468);
or OR2 (N3831, N3828, N2637);
nor NOR3 (N3832, N3829, N2817, N869);
not NOT1 (N3833, N3831);
nand NAND2 (N3834, N3826, N1572);
not NOT1 (N3835, N3821);
and AND3 (N3836, N3824, N3256, N389);
and AND3 (N3837, N3830, N2172, N571);
and AND2 (N3838, N3811, N1833);
nor NOR2 (N3839, N3838, N50);
nor NOR3 (N3840, N3832, N3757, N2041);
nor NOR4 (N3841, N3837, N3245, N1301, N3775);
nor NOR2 (N3842, N3827, N3817);
nand NAND4 (N3843, N3842, N1822, N2682, N1493);
buf BUF1 (N3844, N3834);
xor XOR2 (N3845, N3833, N3123);
nor NOR4 (N3846, N3835, N1305, N205, N2876);
nand NAND3 (N3847, N3841, N534, N1649);
xor XOR2 (N3848, N3823, N88);
nor NOR4 (N3849, N3844, N3711, N3395, N3157);
buf BUF1 (N3850, N3846);
buf BUF1 (N3851, N3850);
and AND4 (N3852, N3848, N2008, N966, N3676);
nor NOR2 (N3853, N3845, N1339);
xor XOR2 (N3854, N3847, N1121);
and AND2 (N3855, N3852, N2892);
buf BUF1 (N3856, N3836);
xor XOR2 (N3857, N3843, N1142);
buf BUF1 (N3858, N3856);
not NOT1 (N3859, N3840);
nand NAND4 (N3860, N3849, N1630, N1639, N2632);
not NOT1 (N3861, N3851);
buf BUF1 (N3862, N3859);
nand NAND3 (N3863, N3860, N2430, N1259);
nand NAND4 (N3864, N3855, N1680, N2474, N2578);
buf BUF1 (N3865, N3857);
nand NAND3 (N3866, N3864, N483, N501);
buf BUF1 (N3867, N3803);
and AND2 (N3868, N3865, N383);
nand NAND2 (N3869, N3863, N710);
or OR3 (N3870, N3862, N2441, N2369);
nor NOR4 (N3871, N3870, N2789, N2042, N298);
buf BUF1 (N3872, N3858);
xor XOR2 (N3873, N3869, N208);
buf BUF1 (N3874, N3866);
xor XOR2 (N3875, N3839, N1389);
or OR2 (N3876, N3875, N3393);
or OR3 (N3877, N3872, N2374, N915);
not NOT1 (N3878, N3871);
nand NAND2 (N3879, N3867, N1422);
and AND2 (N3880, N3876, N3493);
not NOT1 (N3881, N3853);
or OR2 (N3882, N3880, N3337);
nor NOR3 (N3883, N3874, N1610, N276);
xor XOR2 (N3884, N3878, N559);
or OR2 (N3885, N3883, N3142);
buf BUF1 (N3886, N3881);
xor XOR2 (N3887, N3884, N1548);
nand NAND3 (N3888, N3854, N2970, N1853);
buf BUF1 (N3889, N3887);
or OR2 (N3890, N3877, N3345);
and AND2 (N3891, N3873, N869);
not NOT1 (N3892, N3889);
not NOT1 (N3893, N3868);
and AND4 (N3894, N3893, N3106, N3510, N182);
nor NOR4 (N3895, N3891, N3815, N917, N3487);
nor NOR3 (N3896, N3895, N3818, N1791);
nand NAND3 (N3897, N3888, N2841, N465);
and AND2 (N3898, N3861, N2567);
nor NOR4 (N3899, N3898, N2120, N3731, N1705);
and AND3 (N3900, N3896, N2852, N1363);
nor NOR4 (N3901, N3879, N3768, N302, N218);
not NOT1 (N3902, N3892);
or OR4 (N3903, N3902, N1164, N1372, N1404);
and AND4 (N3904, N3900, N2382, N1483, N413);
not NOT1 (N3905, N3882);
nand NAND3 (N3906, N3885, N1336, N1574);
xor XOR2 (N3907, N3906, N1147);
nor NOR3 (N3908, N3903, N134, N784);
nor NOR2 (N3909, N3894, N1817);
or OR3 (N3910, N3901, N2736, N1919);
not NOT1 (N3911, N3910);
buf BUF1 (N3912, N3886);
buf BUF1 (N3913, N3905);
xor XOR2 (N3914, N3908, N3667);
and AND3 (N3915, N3912, N3647, N2737);
xor XOR2 (N3916, N3890, N3367);
nor NOR2 (N3917, N3897, N2065);
and AND3 (N3918, N3915, N2789, N2475);
not NOT1 (N3919, N3918);
and AND3 (N3920, N3914, N3647, N1698);
buf BUF1 (N3921, N3904);
nor NOR3 (N3922, N3913, N3021, N3883);
buf BUF1 (N3923, N3920);
nor NOR4 (N3924, N3911, N2657, N3483, N1859);
and AND2 (N3925, N3907, N3254);
and AND4 (N3926, N3916, N388, N950, N2278);
nand NAND4 (N3927, N3919, N1429, N3766, N271);
xor XOR2 (N3928, N3921, N437);
or OR2 (N3929, N3927, N3851);
and AND4 (N3930, N3924, N2616, N3033, N354);
and AND4 (N3931, N3923, N579, N2655, N1260);
not NOT1 (N3932, N3930);
buf BUF1 (N3933, N3899);
xor XOR2 (N3934, N3909, N1342);
buf BUF1 (N3935, N3925);
not NOT1 (N3936, N3922);
or OR3 (N3937, N3936, N2720, N1795);
or OR3 (N3938, N3932, N2138, N1239);
buf BUF1 (N3939, N3937);
xor XOR2 (N3940, N3917, N2723);
and AND2 (N3941, N3938, N3265);
nor NOR2 (N3942, N3926, N3823);
nand NAND3 (N3943, N3939, N282, N1509);
and AND2 (N3944, N3943, N3094);
nor NOR3 (N3945, N3944, N1125, N2061);
nor NOR2 (N3946, N3928, N1154);
and AND2 (N3947, N3934, N1067);
not NOT1 (N3948, N3935);
and AND2 (N3949, N3941, N286);
and AND2 (N3950, N3929, N890);
and AND3 (N3951, N3945, N3594, N3820);
not NOT1 (N3952, N3933);
nor NOR2 (N3953, N3931, N91);
not NOT1 (N3954, N3949);
and AND4 (N3955, N3940, N772, N3237, N2060);
nand NAND3 (N3956, N3951, N319, N2758);
not NOT1 (N3957, N3953);
nor NOR2 (N3958, N3950, N259);
buf BUF1 (N3959, N3942);
buf BUF1 (N3960, N3956);
xor XOR2 (N3961, N3952, N2298);
nand NAND3 (N3962, N3958, N3383, N3799);
or OR4 (N3963, N3955, N1061, N3583, N1389);
not NOT1 (N3964, N3948);
nor NOR2 (N3965, N3946, N1532);
nand NAND3 (N3966, N3959, N2477, N2546);
or OR2 (N3967, N3966, N1021);
nand NAND4 (N3968, N3957, N116, N3718, N1264);
xor XOR2 (N3969, N3954, N1171);
or OR2 (N3970, N3965, N1763);
not NOT1 (N3971, N3947);
nor NOR3 (N3972, N3964, N1993, N2143);
nor NOR3 (N3973, N3969, N1894, N2073);
nand NAND2 (N3974, N3968, N1780);
nor NOR2 (N3975, N3972, N3224);
and AND4 (N3976, N3974, N1011, N857, N1223);
and AND3 (N3977, N3975, N3341, N968);
or OR3 (N3978, N3971, N2866, N1719);
not NOT1 (N3979, N3967);
or OR2 (N3980, N3973, N3809);
not NOT1 (N3981, N3960);
and AND3 (N3982, N3961, N3123, N595);
buf BUF1 (N3983, N3980);
and AND4 (N3984, N3977, N3943, N3738, N3173);
nor NOR4 (N3985, N3981, N1393, N1017, N124);
xor XOR2 (N3986, N3962, N484);
not NOT1 (N3987, N3984);
nor NOR4 (N3988, N3986, N1752, N822, N771);
buf BUF1 (N3989, N3983);
xor XOR2 (N3990, N3978, N3267);
and AND2 (N3991, N3982, N2160);
buf BUF1 (N3992, N3987);
nor NOR4 (N3993, N3970, N353, N2553, N3312);
and AND2 (N3994, N3990, N1430);
or OR3 (N3995, N3976, N3150, N3699);
nand NAND2 (N3996, N3992, N3521);
nand NAND4 (N3997, N3995, N3402, N1559, N578);
nand NAND4 (N3998, N3997, N1152, N1303, N1990);
nor NOR2 (N3999, N3988, N2747);
nor NOR4 (N4000, N3999, N726, N956, N2520);
buf BUF1 (N4001, N3994);
not NOT1 (N4002, N4001);
buf BUF1 (N4003, N3996);
and AND3 (N4004, N3993, N1835, N2705);
nor NOR2 (N4005, N4000, N1850);
nand NAND3 (N4006, N3963, N2256, N683);
nor NOR2 (N4007, N4002, N2955);
buf BUF1 (N4008, N3998);
not NOT1 (N4009, N4006);
or OR3 (N4010, N3979, N799, N558);
nand NAND2 (N4011, N4003, N3047);
nand NAND2 (N4012, N3985, N1735);
and AND2 (N4013, N4011, N1648);
buf BUF1 (N4014, N4004);
and AND2 (N4015, N4009, N3502);
nor NOR3 (N4016, N4010, N2479, N1470);
not NOT1 (N4017, N4015);
endmodule